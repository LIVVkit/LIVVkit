netcdf dome.diffsmall.10 {
dimensions:
	time = UNLIMITED ; // (11 currently)
	level = 10 ;
	lithoz = 20 ;
	staglevel = 9 ;
	stagwbndlevel = 11 ;
	x0 = 10 ;
	x1 = 11 ;
	y0 = 10 ;
	y1 = 11 ;
variables:
	float time(time) ;
		time:long_name = "Model time" ;
		time:standard_name = "time" ;
		time:units = "year since 1-1-1 0:0:0" ;
		time:calendar = "none" ;
	float level(level) ;
		level:positive = "down" ;
		level:long_name = "sigma layers" ;
		level:standard_name = "land_ice_sigma_coordinate" ;
		level:units = "1" ;
	float lithoz(lithoz) ;
		lithoz:long_name = "vertical coordinate of lithosphere layer" ;
		lithoz:units = "meter" ;
	float staglevel(staglevel) ;
		staglevel:positive = "down" ;
		staglevel:long_name = "stag sigma layers" ;
		staglevel:standard_name = "land_ice_stag_sigma_coordinate" ;
		staglevel:units = "1" ;
	float stagwbndlevel(stagwbndlevel) ;
		stagwbndlevel:positive = "down" ;
		stagwbndlevel:long_name = "stag sigma layers with boundaries" ;
		stagwbndlevel:standard_name = "land_ice_stag_sigma_coordinate_with_bnd" ;
		stagwbndlevel:units = "1" ;
	float x0(x0) ;
		x0:long_name = "Cartesian x-coordinate, velocity grid" ;
		x0:units = "meter" ;
		x0:axis = "X" ;
	float x1(x1) ;
		x1:long_name = "Cartesian x-coordinate" ;
		x1:units = "meter" ;
		x1:axis = "X" ;
	float y0(y0) ;
		y0:long_name = "Cartesian y-coordinate, velocity grid" ;
		y0:units = "meter" ;
		y0:axis = "Y" ;
	float y1(y1) ;
		y1:long_name = "Cartesian y-coordinate" ;
		y1:units = "meter" ;
		y1:axis = "Y" ;
	float tempstag(time, stagwbndlevel, y1, x1) ;
		tempstag:long_name = "ice temperature on staggered vertical levels with boundaries" ;
		tempstag:standard_name = "land_ice_temperature_stag" ;
		tempstag:units = "degree_Celsius" ;
	float thk(time, y1, x1) ;
		thk:scale_factor = 2000. ;
		thk:long_name = "ice thickness" ;
		thk:standard_name = "land_ice_thickness" ;
		thk:units = "meter" ;
	float usurf(time, y1, x1) ;
		usurf:scale_factor = 2000. ;
		usurf:long_name = "ice upper surface elevation" ;
		usurf:standard_name = "surface_altitude" ;
		usurf:units = "meter" ;
	float uvel(time, level, y0, x0) ;
		uvel:scale_factor = 500. ;
		uvel:long_name = "ice velocity in x direction" ;
		uvel:standard_name = "land_ice_x_velocity" ;
		uvel:units = "meter/year" ;
	float velnorm(time, level, y0, x0) ;
		velnorm:scale_factor = 500. ;
		velnorm:long_name = "Horizontal ice velocity magnitude" ;
		velnorm:units = "meter/year" ;
	float vvel(time, level, y0, x0) ;
		vvel:scale_factor = 500. ;
		vvel:long_name = "ice velocity in y direction" ;
		vvel:standard_name = "land_ice_y_velocity" ;
		vvel:units = "meter/year" ;

// global attributes:
		:Conventions = "CF-1.3" ;
		:title = "parabolic dome test case using first-order dynamics" ;
		:institution = "" ;
		:source = "Generated by CISM 2.0" ;
		:history = "2015-05-29 14:19:55.371 : CISM 2.0" ;
		:references = "" ;
		:comment = "created with dome.py" ;
		:configuration = "[DOME-TEST]\n",
			"[grid]\n",
			"upn: 10\n",
			"ewn: 11\n",
			"nsn: 11\n",
			"dew: 6000\n",
			"dns: 6000\n",
			"[time]\n",
			"tstart: 0.\n",
			"tend: 10.\n",
			"dt: 1.\n",
			"dt_diag: 1.\n",
			"idiag: 10\n",
			"jdiag: 10\n",
			"[options]\n",
			"dycore: 2                  # 1 = glam, 2 = glissade\n",
			"flow_law: 2                # 0 = isothermal, 2 = temperature dependent\n",
			"evolution: 3               # 3 = inc. remapping, 4 = FO upwind\n",
			"temperature: 1             # 0 = set column to surf. air temp, 1 = prognostic, 2 = hold at init. values\n",
			"[ho_options]\n",
			"which_ho_babc: 4           # 4 = no-slip at bed\n",
			"which_ho_efvs: 2           # 2 = nonlinear eff. visc. w/ n=3\n",
			"which_ho_sparse: 3         # 1 = SLAP GMRES, 3 = glissade parallel PCG, 4 = Trilinos for linear solver\n",
			"which_ho_nonlinear: 0      # 0 = Picard, 1 = JFNK\n",
			"[parameters]\n",
			"ice_limit: 1.          # min thickness (m) for dynamics\n",
			"[CF default]\n",
			"comment: created with dome.py\n",
			"title: parabolic dome test case using first-order dynamics\n",
			"[CF input]\n",
			"name: dome.nc\n",
			"time: 1\n",
			"[CF output]\n",
			"variables: thk usurf uvel vvel velnorm temp\n",
			"frequency: 1\n",
			"name: dome.base.10.nc\n",
			"" ;
data:

 time = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 level = 0, 0.2533333, 0.4407713, 0.5833333, 0.6942801, 0.7823129, 0.8533334, 
    0.9114583, 0.9596309, 1 ;

 lithoz = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 staglevel = 0.1266667, 0.3470523, 0.5120524, 0.6388067, 0.7382965, 
    0.8178231, 0.8823958, 0.9355446, 0.9798155 ;

 stagwbndlevel = 0, 0.1266667, 0.3470523, 0.5120524, 0.6388067, 0.7382965, 
    0.8178231, 0.8823958, 0.9355446, 0.9798155, 1 ;

 x0 = 3000, 9000, 15000, 21000, 27000, 33000, 39000, 45000, 51000, 57000 ;

 x1 = 0, 6000, 12000, 18000, 24000, 30000, 36000, 42000, 48000, 54000, 60000 ;

 y0 = 3000, 9000, 15000, 21000, 27000, 33000, 39000, 45000, 51000, 57000 ;

 y1 = 0, 6000, 12000, 18000, 24000, 30000, 36000, 42000, 48000, 54000, 60000 ;

 tempstag =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, -15, -15, -15, -15, -15, -15, -15, 0, 0,
  0, 0, 0, -15, -15, -15, -15, -15, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.99997, -14.99983, -14.99967, -14.99983, -14.99997, 0, 0, 0,
  0, 0, -14.99997, -14.99997, -14.99987, -14.99967, -14.99987, -14.99997, 
    -14.99997, 0, 0,
  0, -14.99997, -14.99997, -14.99997, -14.99996, -14.99995, -14.99996, 
    -14.99997, -14.99997, -14.99997, 0,
  0, -14.99983, -14.99987, -14.99996, -14.99998, -14.99999, -14.99998, 
    -14.99996, -14.99987, -14.99983, 0,
  0, -14.99967, -14.99967, -14.99995, -14.99999, -15, -14.99999, -14.99995, 
    -14.99967, -14.99967, 0,
  0, -14.99983, -14.99987, -14.99996, -14.99998, -14.99999, -14.99998, 
    -14.99996, -14.99987, -14.99983, 0,
  0, -14.99997, -14.99997, -14.99997, -14.99996, -14.99995, -14.99996, 
    -14.99997, -14.99997, -14.99997, 0,
  0, 0, -14.99997, -14.99997, -14.99987, -14.99967, -14.99987, -14.99997, 
    -14.99997, 0, 0,
  0, 0, 0, -14.99997, -14.99983, -14.99967, -14.99983, -14.99997, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.99993, -14.99973, -14.99956, -14.99973, -14.99993, 0, 0, 0,
  0, 0, -14.99994, -14.99992, -14.99975, -14.9995, -14.99975, -14.99992, 
    -14.99994, 0, 0,
  0, -14.99993, -14.99992, -14.99993, -14.99993, -14.99993, -14.99993, 
    -14.99993, -14.99992, -14.99993, 0,
  0, -14.99973, -14.99975, -14.99993, -14.99998, -14.99999, -14.99998, 
    -14.99993, -14.99975, -14.99973, 0,
  0, -14.99956, -14.9995, -14.99993, -14.99999, -15, -14.99999, -14.99993, 
    -14.9995, -14.99956, 0,
  0, -14.99973, -14.99975, -14.99993, -14.99998, -14.99999, -14.99998, 
    -14.99993, -14.99975, -14.99973, 0,
  0, -14.99993, -14.99992, -14.99993, -14.99993, -14.99993, -14.99993, 
    -14.99993, -14.99992, -14.99993, 0,
  0, 0, -14.99994, -14.99992, -14.99975, -14.9995, -14.99975, -14.99992, 
    -14.99994, 0, 0,
  0, 0, 0, -14.99993, -14.99973, -14.99956, -14.99973, -14.99993, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.99987, -14.99955, -14.99936, -14.99955, -14.99987, 0, 0, 0,
  0, 0, -14.99991, -14.99974, -14.99935, -14.99895, -14.99935, -14.99974, 
    -14.99991, 0, 0,
  0, -14.99987, -14.99974, -14.99976, -14.99985, -14.99987, -14.99985, 
    -14.99976, -14.99974, -14.99987, 0,
  0, -14.99955, -14.99935, -14.99985, -14.99997, -14.99999, -14.99997, 
    -14.99985, -14.99935, -14.99955, 0,
  0, -14.99936, -14.99895, -14.99987, -14.99999, -15, -14.99999, -14.99987, 
    -14.99895, -14.99936, 0,
  0, -14.99955, -14.99935, -14.99985, -14.99997, -14.99999, -14.99997, 
    -14.99985, -14.99935, -14.99955, 0,
  0, -14.99987, -14.99974, -14.99976, -14.99985, -14.99987, -14.99985, 
    -14.99976, -14.99974, -14.99987, 0,
  0, 0, -14.99991, -14.99974, -14.99935, -14.99895, -14.99935, -14.99974, 
    -14.99991, 0, 0,
  0, 0, 0, -14.99987, -14.99955, -14.99936, -14.99955, -14.99987, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.99969, -14.99916, -14.99895, -14.99916, -14.99969, 0, 0, 0,
  0, 0, -14.99985, -14.99941, -14.99856, -14.99786, -14.99856, -14.99941, 
    -14.99985, 0, 0,
  0, -14.99969, -14.99941, -14.99944, -14.99971, -14.99978, -14.99971, 
    -14.99944, -14.99941, -14.99969, 0,
  0, -14.99916, -14.99856, -14.99971, -14.99994, -14.99998, -14.99994, 
    -14.99971, -14.99856, -14.99916, 0,
  0, -14.99895, -14.99786, -14.99978, -14.99998, -15, -14.99998, -14.99978, 
    -14.99786, -14.99895, 0,
  0, -14.99916, -14.99856, -14.99971, -14.99994, -14.99998, -14.99994, 
    -14.99971, -14.99856, -14.99916, 0,
  0, -14.99969, -14.99941, -14.99944, -14.99971, -14.99978, -14.99971, 
    -14.99944, -14.99941, -14.99969, 0,
  0, 0, -14.99985, -14.99941, -14.99856, -14.99786, -14.99856, -14.99941, 
    -14.99985, 0, 0,
  0, 0, 0, -14.99969, -14.99916, -14.99895, -14.99916, -14.99969, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.99942, -14.99834, -14.99806, -14.99834, -14.99942, 0, 0, 0,
  0, 0, -14.9997, -14.99897, -14.99744, -14.99628, -14.99744, -14.99897, 
    -14.9997, 0, 0,
  0, -14.99942, -14.99897, -14.999, -14.99951, -14.99966, -14.99951, -14.999, 
    -14.99897, -14.99942, 0,
  0, -14.99834, -14.99744, -14.99951, -14.99991, -14.99997, -14.99991, 
    -14.99951, -14.99744, -14.99834, 0,
  0, -14.99806, -14.99628, -14.99966, -14.99997, -15, -14.99997, -14.99966, 
    -14.99628, -14.99806, 0,
  0, -14.99834, -14.99744, -14.99951, -14.99991, -14.99997, -14.99991, 
    -14.99951, -14.99744, -14.99834, 0,
  0, -14.99942, -14.99897, -14.999, -14.99951, -14.99966, -14.99951, -14.999, 
    -14.99897, -14.99942, 0,
  0, 0, -14.9997, -14.99897, -14.99744, -14.99628, -14.99744, -14.99897, 
    -14.9997, 0, 0,
  0, 0, 0, -14.99942, -14.99834, -14.99806, -14.99834, -14.99942, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.99917, -14.99761, -14.99724, -14.99761, -14.99917, 0, 0, 0,
  0, 0, -14.99957, -14.99834, -14.99611, -14.99438, -14.99611, -14.99834, 
    -14.99957, 0, 0,
  0, -14.99917, -14.99834, -14.99847, -14.99927, -14.99951, -14.99927, 
    -14.99847, -14.99834, -14.99917, 0,
  0, -14.99761, -14.99611, -14.99927, -14.99988, -14.99996, -14.99988, 
    -14.99927, -14.99611, -14.99761, 0,
  0, -14.99724, -14.99438, -14.99951, -14.99996, -15, -14.99996, -14.99951, 
    -14.99438, -14.99724, 0,
  0, -14.99761, -14.99611, -14.99927, -14.99988, -14.99996, -14.99988, 
    -14.99927, -14.99611, -14.99761, 0,
  0, -14.99917, -14.99834, -14.99847, -14.99927, -14.99951, -14.99927, 
    -14.99847, -14.99834, -14.99917, 0,
  0, 0, -14.99957, -14.99834, -14.99611, -14.99438, -14.99611, -14.99834, 
    -14.99957, 0, 0,
  0, 0, 0, -14.99917, -14.99761, -14.99724, -14.99761, -14.99917, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.99876, -14.99652, -14.996, -14.99652, -14.99876, 0, 0, 0,
  0, 0, -14.99936, -14.99652, -14.99445, -14.99215, -14.99445, -14.99652, 
    -14.99936, 0, 0,
  0, -14.99876, -14.99652, -14.9978, -14.99897, -14.9993, -14.99897, 
    -14.9978, -14.99652, -14.99876, 0,
  0, -14.99652, -14.99445, -14.99897, -14.99981, -14.99993, -14.99981, 
    -14.99897, -14.99445, -14.99652, 0,
  0, -14.996, -14.99215, -14.9993, -14.99993, -14.99998, -14.99993, -14.9993, 
    -14.99215, -14.996, 0,
  0, -14.99652, -14.99445, -14.99897, -14.99981, -14.99993, -14.99981, 
    -14.99897, -14.99445, -14.99652, 0,
  0, -14.99876, -14.99652, -14.9978, -14.99897, -14.9993, -14.99897, 
    -14.9978, -14.99652, -14.99876, 0,
  0, 0, -14.99936, -14.99652, -14.99445, -14.99215, -14.99445, -14.99652, 
    -14.99936, 0, 0,
  0, 0, 0, -14.99876, -14.99652, -14.996, -14.99652, -14.99876, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.99789, -14.99477, -14.99405, -14.99477, -14.99789, 0, 0, 0,
  0, 0, -14.99877, -14.98636, -14.98925, -14.987, -14.98925, -14.98636, 
    -14.99877, 0, 0,
  0, -14.99789, -14.98636, -14.99474, -14.99713, -14.99775, -14.99713, 
    -14.99474, -14.98636, -14.99789, 0,
  0, -14.99477, -14.98925, -14.99713, -14.99865, -14.99891, -14.99865, 
    -14.99713, -14.98925, -14.99477, 0,
  0, -14.99405, -14.987, -14.99775, -14.99891, -14.99907, -14.99891, 
    -14.99775, -14.987, -14.99405, 0,
  0, -14.99477, -14.98925, -14.99713, -14.99865, -14.99891, -14.99865, 
    -14.99713, -14.98925, -14.99477, 0,
  0, -14.99789, -14.98636, -14.99474, -14.99713, -14.99775, -14.99713, 
    -14.99474, -14.98636, -14.99789, 0,
  0, 0, -14.99877, -14.98636, -14.98925, -14.987, -14.98925, -14.98636, 
    -14.99877, 0, 0,
  0, 0, 0, -14.99789, -14.99477, -14.99405, -14.99477, -14.99789, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -14.9868, -14.98577, -14.98567, -14.98577, -14.9868, 0, 0, 0,
  0, 0, -14.98722, -14.93203, -14.94519, -14.94489, -14.94519, -14.93203, 
    -14.98722, 0, 0,
  0, -14.9868, -14.93203, -14.95609, -14.96362, -14.96558, -14.96362, 
    -14.95609, -14.93203, -14.9868, 0,
  0, -14.98577, -14.94519, -14.96362, -14.96872, -14.96992, -14.96872, 
    -14.96362, -14.94519, -14.98577, 0,
  0, -14.98567, -14.94489, -14.96558, -14.96992, -14.97093, -14.96992, 
    -14.96558, -14.94489, -14.98567, 0,
  0, -14.98577, -14.94519, -14.96362, -14.96872, -14.96992, -14.96872, 
    -14.96362, -14.94519, -14.98577, 0,
  0, -14.9868, -14.93203, -14.95609, -14.96362, -14.96558, -14.96362, 
    -14.95609, -14.93203, -14.9868, 0,
  0, 0, -14.98722, -14.93203, -14.94519, -14.94489, -14.94519, -14.93203, 
    -14.98722, 0, 0,
  0, 0, 0, -14.9868, -14.98577, -14.98567, -14.98577, -14.9868, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -14.80461, -14.74738, -14.72864, -14.74738, -14.80461, -15, 
    -15, -15,
  -15, -15, -14.80461, -14.72285, -14.68559, -14.67413, -14.68559, -14.72285, 
    -14.80461, -15, -15,
  -15, -15, -14.74738, -14.68559, -14.65216, -14.64153, -14.65216, -14.68559, 
    -14.74738, -15, -15,
  -15, -15, -14.72864, -14.67413, -14.64153, -14.6311, -14.64153, -14.67413, 
    -14.72864, -15, -15,
  -15, -15, -14.74738, -14.68559, -14.65216, -14.64153, -14.65216, -14.68559, 
    -14.74738, -15, -15,
  -15, -15, -14.80461, -14.72285, -14.68559, -14.67413, -14.68559, -14.72285, 
    -14.80461, -15, -15,
  -15, -15, -15, -14.80461, -14.74738, -14.72864, -14.74738, -14.80461, -15, 
    -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99997, -14.99996, -14.9974, -14.99996, -14.99997, -15, 0, 0,
  0, -15, -14.99999, -14.99994, -14.99985, -14.99966, -14.99985, -14.99994, 
    -14.99999, -15, 0,
  0, -14.99997, -14.99994, -14.99995, -14.99992, -14.99991, -14.99992, 
    -14.99995, -14.99994, -14.99997, 0,
  0, -14.99996, -14.99985, -14.99992, -14.99996, -14.99999, -14.99996, 
    -14.99992, -14.99985, -14.99996, 0,
  0, -14.9974, -14.99966, -14.99991, -14.99999, -15, -14.99999, -14.99991, 
    -14.99966, -14.9974, 0,
  0, -14.99996, -14.99985, -14.99992, -14.99996, -14.99999, -14.99996, 
    -14.99992, -14.99985, -14.99996, 0,
  0, -14.99997, -14.99994, -14.99995, -14.99992, -14.99991, -14.99992, 
    -14.99995, -14.99994, -14.99997, 0,
  0, -15, -14.99999, -14.99994, -14.99985, -14.99966, -14.99985, -14.99994, 
    -14.99999, -15, 0,
  0, 0, -15, -14.99997, -14.99996, -14.9974, -14.99996, -14.99997, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99992, -14.99991, -14.99326, -14.99991, -14.99992, -15, 0, 0,
  0, -15, -14.99996, -14.99983, -14.99966, -14.99941, -14.99966, -14.99983, 
    -14.99996, -15, 0,
  0, -14.99992, -14.99983, -14.99985, -14.99986, -14.99986, -14.99986, 
    -14.99985, -14.99983, -14.99992, 0,
  0, -14.99991, -14.99966, -14.99986, -14.99995, -14.99998, -14.99995, 
    -14.99986, -14.99966, -14.99991, 0,
  0, -14.99326, -14.99941, -14.99986, -14.99998, -15, -14.99998, -14.99986, 
    -14.99941, -14.99326, 0,
  0, -14.99991, -14.99966, -14.99986, -14.99995, -14.99998, -14.99995, 
    -14.99986, -14.99966, -14.99991, 0,
  0, -14.99992, -14.99983, -14.99985, -14.99986, -14.99986, -14.99986, 
    -14.99985, -14.99983, -14.99992, 0,
  0, -15, -14.99996, -14.99983, -14.99966, -14.99941, -14.99966, -14.99983, 
    -14.99996, -15, 0,
  0, 0, -15, -14.99992, -14.99991, -14.99326, -14.99991, -14.99992, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99979, -14.99976, -14.98982, -14.99976, -14.99979, -15, 0, 0,
  0, -15, -14.99988, -14.99946, -14.99901, -14.99864, -14.99901, -14.99946, 
    -14.99988, -15, 0,
  0, -14.99979, -14.99946, -14.99952, -14.99971, -14.99976, -14.99971, 
    -14.99952, -14.99946, -14.99979, 0,
  0, -14.99976, -14.99901, -14.99971, -14.99993, -14.99997, -14.99993, 
    -14.99971, -14.99901, -14.99976, 0,
  0, -14.98982, -14.99864, -14.99976, -14.99997, -15, -14.99997, -14.99976, 
    -14.99864, -14.98982, 0,
  0, -14.99976, -14.99901, -14.99971, -14.99993, -14.99997, -14.99993, 
    -14.99971, -14.99901, -14.99976, 0,
  0, -14.99979, -14.99946, -14.99952, -14.99971, -14.99976, -14.99971, 
    -14.99952, -14.99946, -14.99979, 0,
  0, -15, -14.99988, -14.99946, -14.99901, -14.99864, -14.99901, -14.99946, 
    -14.99988, -15, 0,
  0, 0, -15, -14.99979, -14.99976, -14.98982, -14.99976, -14.99979, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.9996, -14.99951, -14.9867, -14.99951, -14.9996, -15, 0, 0,
  0, -15, -14.99977, -14.9988, -14.99774, -14.99712, -14.99774, -14.9988, 
    -14.99977, -15, 0,
  0, -14.9996, -14.9988, -14.99889, -14.99942, -14.99957, -14.99942, 
    -14.99889, -14.9988, -14.9996, 0,
  0, -14.99951, -14.99774, -14.99942, -14.99989, -14.99996, -14.99989, 
    -14.99942, -14.99774, -14.99951, 0,
  0, -14.9867, -14.99712, -14.99957, -14.99996, -15, -14.99996, -14.99957, 
    -14.99712, -14.9867, 0,
  0, -14.99951, -14.99774, -14.99942, -14.99989, -14.99996, -14.99989, 
    -14.99942, -14.99774, -14.99951, 0,
  0, -14.9996, -14.9988, -14.99889, -14.99942, -14.99957, -14.99942, 
    -14.99889, -14.9988, -14.9996, 0,
  0, -15, -14.99977, -14.9988, -14.99774, -14.99712, -14.99774, -14.9988, 
    -14.99977, -15, 0,
  0, 0, -15, -14.9996, -14.99951, -14.9867, -14.99951, -14.9996, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99933, -14.99921, -14.98397, -14.99921, -14.99933, -15, 0, 0,
  0, -15, -14.99962, -14.99788, -14.99597, -14.99497, -14.99597, -14.99788, 
    -14.99962, -15, 0,
  0, -14.99933, -14.99788, -14.998, -14.99902, -14.99931, -14.99902, -14.998, 
    -14.99788, -14.99933, 0,
  0, -14.99921, -14.99597, -14.99902, -14.99983, -14.99995, -14.99983, 
    -14.99902, -14.99597, -14.99921, 0,
  0, -14.98397, -14.99497, -14.99931, -14.99995, -15, -14.99995, -14.99931, 
    -14.99497, -14.98397, 0,
  0, -14.99921, -14.99597, -14.99902, -14.99983, -14.99995, -14.99983, 
    -14.99902, -14.99597, -14.99921, 0,
  0, -14.99933, -14.99788, -14.998, -14.99902, -14.99931, -14.99902, -14.998, 
    -14.99788, -14.99933, 0,
  0, -15, -14.99962, -14.99788, -14.99597, -14.99497, -14.99597, -14.99788, 
    -14.99962, -15, 0,
  0, 0, -15, -14.99933, -14.99921, -14.98397, -14.99921, -14.99933, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99898, -14.99894, -14.9816, -14.99894, -14.99898, -15, 0, 0,
  0, -15, -14.99942, -14.99635, -14.99384, -14.99237, -14.99384, -14.99635, 
    -14.99942, -15, 0,
  0, -14.99898, -14.99635, -14.99694, -14.99853, -14.99899, -14.99853, 
    -14.99694, -14.99635, -14.99898, 0,
  0, -14.99894, -14.99384, -14.99853, -14.99975, -14.99993, -14.99975, 
    -14.99853, -14.99384, -14.99894, 0,
  0, -14.9816, -14.99237, -14.99899, -14.99993, -15, -14.99993, -14.99899, 
    -14.99237, -14.9816, 0,
  0, -14.99894, -14.99384, -14.99853, -14.99975, -14.99993, -14.99975, 
    -14.99853, -14.99384, -14.99894, 0,
  0, -14.99898, -14.99635, -14.99694, -14.99853, -14.99899, -14.99853, 
    -14.99694, -14.99635, -14.99898, 0,
  0, -15, -14.99942, -14.99635, -14.99384, -14.99237, -14.99384, -14.99635, 
    -14.99942, -15, 0,
  0, 0, -15, -14.99898, -14.99894, -14.9816, -14.99894, -14.99898, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99837, -14.99873, -14.9795, -14.99873, -14.99837, -15, 0, 0,
  0, -15, -14.99885, -14.99107, -14.99075, -14.98899, -14.99075, -14.99107, 
    -14.99885, -15, 0,
  0, -14.99837, -14.99107, -14.99539, -14.99782, -14.99848, -14.99782, 
    -14.99539, -14.99107, -14.99837, 0,
  0, -14.99873, -14.99075, -14.99782, -14.99956, -14.99981, -14.99956, 
    -14.99782, -14.99075, -14.99873, 0,
  0, -14.9795, -14.98899, -14.99848, -14.99981, -14.99992, -14.99981, 
    -14.99848, -14.98899, -14.9795, 0,
  0, -14.99873, -14.99075, -14.99782, -14.99956, -14.99981, -14.99956, 
    -14.99782, -14.99075, -14.99873, 0,
  0, -14.99837, -14.99107, -14.99539, -14.99782, -14.99848, -14.99782, 
    -14.99539, -14.99107, -14.99837, 0,
  0, -15, -14.99885, -14.99107, -14.99075, -14.98899, -14.99075, -14.99107, 
    -14.99885, -15, 0,
  0, 0, -15, -14.99837, -14.99873, -14.9795, -14.99873, -14.99837, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99565, -14.99829, -14.97757, -14.99829, -14.99565, -15, 0, 0,
  0, -15, -14.99588, -14.96654, -14.97839, -14.97788, -14.97839, -14.96654, 
    -14.99588, -15, 0,
  0, -14.99565, -14.96654, -14.98736, -14.99281, -14.99416, -14.99281, 
    -14.98736, -14.96654, -14.99565, 0,
  0, -14.99829, -14.97839, -14.99281, -14.99629, -14.99691, -14.99629, 
    -14.99281, -14.97839, -14.99829, 0,
  0, -14.97757, -14.97788, -14.99416, -14.99691, -14.99729, -14.99691, 
    -14.99416, -14.97788, -14.97757, 0,
  0, -14.99829, -14.97839, -14.99281, -14.99629, -14.99691, -14.99629, 
    -14.99281, -14.97839, -14.99829, 0,
  0, -14.99565, -14.96654, -14.98736, -14.99281, -14.99416, -14.99281, 
    -14.98736, -14.96654, -14.99565, 0,
  0, -15, -14.99588, -14.96654, -14.97839, -14.97788, -14.97839, -14.96654, 
    -14.99588, -15, 0,
  0, 0, -15, -14.99565, -14.99829, -14.97757, -14.99829, -14.99565, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.98927, -14.99734, -14.97501, -14.99734, -14.98927, -15, 0, 0,
  0, -15, -14.99051, -14.87481, -14.89819, -14.90092, -14.89819, -14.87481, 
    -14.99051, -15, 0,
  0, -14.98927, -14.87481, -14.91507, -14.92902, -14.93266, -14.92902, 
    -14.91507, -14.87481, -14.98927, 0,
  0, -14.99734, -14.89819, -14.92902, -14.93872, -14.94101, -14.93872, 
    -14.92902, -14.89819, -14.99734, 0,
  0, -14.97501, -14.90092, -14.93266, -14.94101, -14.94291, -14.94101, 
    -14.93266, -14.90092, -14.97501, 0,
  0, -14.99734, -14.89819, -14.92902, -14.93872, -14.94101, -14.93872, 
    -14.92902, -14.89819, -14.99734, 0,
  0, -14.98927, -14.87481, -14.91507, -14.92902, -14.93266, -14.92902, 
    -14.91507, -14.87481, -14.98927, 0,
  0, -15, -14.99051, -14.87481, -14.89819, -14.90092, -14.89819, -14.87481, 
    -14.99051, -15, 0,
  0, 0, -15, -14.98927, -14.99734, -14.97501, -14.99734, -14.98927, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -14.97554, -15, -15, -15, -15, -15,
  -15, -15, -15, -14.74725, -14.70049, -14.68504, -14.70049, -14.74725, -15, 
    -15, -15,
  -15, -15, -14.74725, -14.68189, -14.65114, -14.6414, -14.65114, -14.68189, 
    -14.74725, -15, -15,
  -15, -15, -14.70049, -14.65114, -14.62228, -14.61267, -14.62228, -14.65114, 
    -14.70049, -15, -15,
  -15, -14.97554, -14.68504, -14.6414, -14.61267, -14.6031, -14.61267, 
    -14.6414, -14.68504, -14.97554, -15,
  -15, -15, -14.70049, -14.65114, -14.62228, -14.61267, -14.62228, -14.65114, 
    -14.70049, -15, -15,
  -15, -15, -14.74725, -14.68189, -14.65114, -14.6414, -14.65114, -14.68189, 
    -14.74725, -15, -15,
  -15, -15, -15, -14.74725, -14.70049, -14.68504, -14.70049, -14.74725, -15, 
    -15, -15,
  -15, -15, -15, -15, -15, -14.97554, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99997, -14.99997, -14.99677, -14.99997, -14.99997, -15, 0, 0,
  0, -15, -14.99998, -14.99992, -14.99984, -14.99965, -14.99984, -14.99992, 
    -14.99998, -15, 0,
  0, -14.99997, -14.99992, -14.99992, -14.99988, -14.99986, -14.99988, 
    -14.99992, -14.99992, -14.99997, 0,
  0, -14.99997, -14.99984, -14.99988, -14.99995, -14.99998, -14.99995, 
    -14.99988, -14.99984, -14.99997, 0,
  0, -14.99677, -14.99965, -14.99986, -14.99998, -15, -14.99998, -14.99986, 
    -14.99965, -14.99677, 0,
  0, -14.99997, -14.99984, -14.99988, -14.99995, -14.99998, -14.99995, 
    -14.99988, -14.99984, -14.99997, 0,
  0, -14.99997, -14.99992, -14.99992, -14.99988, -14.99986, -14.99988, 
    -14.99992, -14.99992, -14.99997, 0,
  0, -15, -14.99998, -14.99992, -14.99984, -14.99965, -14.99984, -14.99992, 
    -14.99998, -15, 0,
  0, 0, -15, -14.99997, -14.99997, -14.99677, -14.99997, -14.99997, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99991, -14.99991, -14.99152, -14.99991, -14.99991, -15, 0, 0,
  0, -15, -14.99994, -14.99974, -14.99957, -14.99933, -14.99957, -14.99974, 
    -14.99994, -15, 0,
  0, -14.99991, -14.99974, -14.99978, -14.9998, -14.9998, -14.9998, 
    -14.99978, -14.99974, -14.99991, 0,
  0, -14.99991, -14.99957, -14.9998, -14.99993, -14.99997, -14.99993, 
    -14.9998, -14.99957, -14.99991, 0,
  0, -14.99152, -14.99933, -14.9998, -14.99997, -15, -14.99997, -14.9998, 
    -14.99933, -14.99152, 0,
  0, -14.99991, -14.99957, -14.9998, -14.99993, -14.99997, -14.99993, 
    -14.9998, -14.99957, -14.99991, 0,
  0, -14.99991, -14.99974, -14.99978, -14.9998, -14.9998, -14.9998, 
    -14.99978, -14.99974, -14.99991, 0,
  0, -15, -14.99994, -14.99974, -14.99957, -14.99933, -14.99957, -14.99974, 
    -14.99994, -15, 0,
  0, 0, -15, -14.99991, -14.99991, -14.99152, -14.99991, -14.99991, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99976, -14.99974, -14.98722, -14.99974, -14.99976, -15, 0, 0,
  0, -15, -14.99985, -14.99918, -14.99866, -14.99833, -14.99866, -14.99918, 
    -14.99985, -15, 0,
  0, -14.99976, -14.99918, -14.99928, -14.99957, -14.99965, -14.99957, 
    -14.99928, -14.99918, -14.99976, 0,
  0, -14.99974, -14.99866, -14.99957, -14.99989, -14.99996, -14.99989, 
    -14.99957, -14.99866, -14.99974, 0,
  0, -14.98722, -14.99833, -14.99965, -14.99996, -15, -14.99996, -14.99965, 
    -14.99833, -14.98722, 0,
  0, -14.99974, -14.99866, -14.99957, -14.99989, -14.99996, -14.99989, 
    -14.99957, -14.99866, -14.99974, 0,
  0, -14.99976, -14.99918, -14.99928, -14.99957, -14.99965, -14.99957, 
    -14.99928, -14.99918, -14.99976, 0,
  0, -15, -14.99985, -14.99918, -14.99866, -14.99833, -14.99866, -14.99918, 
    -14.99985, -15, 0,
  0, 0, -15, -14.99976, -14.99974, -14.98722, -14.99974, -14.99976, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99954, -14.99946, -14.98338, -14.99946, -14.99954, -15, 0, 0,
  0, -15, -14.9997, -14.99818, -14.99692, -14.99639, -14.99692, -14.99818, 
    -14.9997, -15, 0,
  0, -14.99954, -14.99818, -14.99833, -14.99913, -14.99936, -14.99913, 
    -14.99833, -14.99818, -14.99954, 0,
  0, -14.99946, -14.99692, -14.99913, -14.99983, -14.99994, -14.99983, 
    -14.99913, -14.99692, -14.99946, 0,
  0, -14.98338, -14.99639, -14.99936, -14.99994, -15, -14.99994, -14.99936, 
    -14.99639, -14.98338, 0,
  0, -14.99946, -14.99692, -14.99913, -14.99983, -14.99994, -14.99983, 
    -14.99913, -14.99692, -14.99946, 0,
  0, -14.99954, -14.99818, -14.99833, -14.99913, -14.99936, -14.99913, 
    -14.99833, -14.99818, -14.99954, 0,
  0, -15, -14.9997, -14.99818, -14.99692, -14.99639, -14.99692, -14.99818, 
    -14.9997, -15, 0,
  0, 0, -15, -14.99954, -14.99946, -14.98338, -14.99946, -14.99954, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99924, -14.99913, -14.98011, -14.99913, -14.99924, -15, 0, 0,
  0, -15, -14.99952, -14.99672, -14.9945, -14.99365, -14.9945, -14.99672, 
    -14.99952, -15, 0,
  0, -14.99924, -14.99672, -14.997, -14.99853, -14.99896, -14.99853, -14.997, 
    -14.99672, -14.99924, 0,
  0, -14.99913, -14.9945, -14.99853, -14.99974, -14.99992, -14.99974, 
    -14.99853, -14.9945, -14.99913, 0,
  0, -14.98011, -14.99365, -14.99896, -14.99992, -15, -14.99992, -14.99896, 
    -14.99365, -14.98011, 0,
  0, -14.99913, -14.9945, -14.99853, -14.99974, -14.99992, -14.99974, 
    -14.99853, -14.9945, -14.99913, 0,
  0, -14.99924, -14.99672, -14.997, -14.99853, -14.99896, -14.99853, -14.997, 
    -14.99672, -14.99924, 0,
  0, -15, -14.99952, -14.99672, -14.9945, -14.99365, -14.9945, -14.99672, 
    -14.99952, -15, 0,
  0, 0, -15, -14.99924, -14.99913, -14.98011, -14.99913, -14.99924, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99882, -14.99885, -14.97731, -14.99885, -14.99882, -15, 0, 0,
  0, -15, -14.99918, -14.99392, -14.99152, -14.99033, -14.99152, -14.99392, 
    -14.99918, -15, 0,
  0, -14.99882, -14.99392, -14.99539, -14.99779, -14.99846, -14.99779, 
    -14.99539, -14.99392, -14.99882, 0,
  0, -14.99885, -14.99152, -14.99779, -14.99963, -14.99989, -14.99963, 
    -14.99779, -14.99152, -14.99885, 0,
  0, -14.97731, -14.99033, -14.99846, -14.99989, -15, -14.99989, -14.99846, 
    -14.99033, -14.97731, 0,
  0, -14.99885, -14.99152, -14.99779, -14.99963, -14.99989, -14.99963, 
    -14.99779, -14.99152, -14.99885, 0,
  0, -14.99882, -14.99392, -14.99539, -14.99779, -14.99846, -14.99779, 
    -14.99539, -14.99392, -14.99882, 0,
  0, -15, -14.99918, -14.99392, -14.99152, -14.99033, -14.99152, -14.99392, 
    -14.99918, -15, 0,
  0, 0, -15, -14.99882, -14.99885, -14.97731, -14.99885, -14.99882, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99771, -14.9986, -14.97481, -14.9986, -14.99771, -15, 0, 0,
  0, -15, -14.99799, -14.98371, -14.98655, -14.98546, -14.98655, -14.98371, 
    -14.99799, -15, 0,
  0, -14.99771, -14.98371, -14.99272, -14.99654, -14.99755, -14.99654, 
    -14.99272, -14.98371, -14.99771, 0,
  0, -14.9986, -14.98655, -14.99654, -14.99924, -14.99963, -14.99924, 
    -14.99654, -14.98655, -14.9986, 0,
  0, -14.97481, -14.98546, -14.99755, -14.99963, -14.9998, -14.99963, 
    -14.99755, -14.98546, -14.97481, 0,
  0, -14.9986, -14.98655, -14.99654, -14.99924, -14.99963, -14.99924, 
    -14.99654, -14.98655, -14.9986, 0,
  0, -14.99771, -14.98371, -14.99272, -14.99654, -14.99755, -14.99654, 
    -14.99272, -14.98371, -14.99771, 0,
  0, -15, -14.99799, -14.98371, -14.98655, -14.98546, -14.98655, -14.98371, 
    -14.99799, -15, 0,
  0, 0, -15, -14.99771, -14.9986, -14.97481, -14.9986, -14.99771, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99448, -14.99793, -14.97238, -14.99793, -14.99448, -15, 0, 0,
  0, -15, -14.99473, -14.94353, -14.96525, -14.96679, -14.96525, -14.94353, 
    -14.99473, -15, 0,
  0, -14.99448, -14.94353, -14.97825, -14.98727, -14.98946, -14.98727, 
    -14.97825, -14.94353, -14.99448, 0,
  0, -14.99793, -14.96525, -14.98727, -14.99301, -14.99406, -14.99301, 
    -14.98727, -14.96525, -14.99793, 0,
  0, -14.97238, -14.96679, -14.98946, -14.99406, -14.99476, -14.99406, 
    -14.98946, -14.96679, -14.97238, 0,
  0, -14.99793, -14.96525, -14.98727, -14.99301, -14.99406, -14.99301, 
    -14.98727, -14.96525, -14.99793, 0,
  0, -14.99448, -14.94353, -14.97825, -14.98727, -14.98946, -14.98727, 
    -14.97825, -14.94353, -14.99448, 0,
  0, -15, -14.99473, -14.94353, -14.96525, -14.96679, -14.96525, -14.94353, 
    -14.99473, -15, 0,
  0, 0, -15, -14.99448, -14.99793, -14.97238, -14.99793, -14.99448, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99158, -14.99707, -14.96953, -14.99707, -14.99158, -15, 0, 0,
  0, -15, -14.99216, -14.82525, -14.85481, -14.85995, -14.85481, -14.82525, 
    -14.99216, -15, 0,
  0, -14.99158, -14.82525, -14.87658, -14.89606, -14.90119, -14.89606, 
    -14.87658, -14.82525, -14.99158, 0,
  0, -14.99707, -14.85481, -14.89606, -14.90991, -14.91318, -14.90991, 
    -14.89606, -14.85481, -14.99707, 0,
  0, -14.96953, -14.85995, -14.90119, -14.91318, -14.9159, -14.91318, 
    -14.90119, -14.85995, -14.96953, 0,
  0, -14.99707, -14.85481, -14.89606, -14.90991, -14.91318, -14.90991, 
    -14.89606, -14.85481, -14.99707, 0,
  0, -14.99158, -14.82525, -14.87658, -14.89606, -14.90119, -14.89606, 
    -14.87658, -14.82525, -14.99158, 0,
  0, -15, -14.99216, -14.82525, -14.85481, -14.85995, -14.85481, -14.82525, 
    -14.99216, -15, 0,
  0, 0, -15, -14.99158, -14.99707, -14.96953, -14.99707, -14.99158, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -14.97029, -15, -15, -15, -15, -15,
  -15, -15, -15, -14.69756, -14.65708, -14.64403, -14.65708, -14.69756, -15, 
    -15, -15,
  -15, -15, -14.69756, -14.64345, -14.61835, -14.61014, -14.61835, -14.64345, 
    -14.69756, -15, -15,
  -15, -15, -14.65708, -14.61835, -14.59358, -14.5849, -14.59358, -14.61835, 
    -14.65708, -15, -15,
  -15, -14.97029, -14.64403, -14.61014, -14.5849, -14.57609, -14.5849, 
    -14.61014, -14.64403, -14.97029, -15,
  -15, -15, -14.65708, -14.61835, -14.59358, -14.5849, -14.59358, -14.61835, 
    -14.65708, -15, -15,
  -15, -15, -14.69756, -14.64345, -14.61835, -14.61014, -14.61835, -14.64345, 
    -14.69756, -15, -15,
  -15, -15, -15, -14.69756, -14.65708, -14.64403, -14.65708, -14.69756, -15, 
    -15, -15,
  -15, -15, -15, -15, -15, -14.97029, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99999, -14.99711, -14.99581, -14.99711, -14.99999, -15, 0, 0,
  0, -15, -14.99998, -14.99988, -14.99981, -14.99963, -14.99981, -14.99988, 
    -14.99998, -15, 0,
  0, -14.99999, -14.99988, -14.99989, -14.99984, -14.99983, -14.99984, 
    -14.99989, -14.99988, -14.99999, 0,
  0, -14.99711, -14.99981, -14.99984, -14.99993, -14.99997, -14.99993, 
    -14.99984, -14.99981, -14.99711, 0,
  0, -14.99581, -14.99963, -14.99983, -14.99997, -15, -14.99997, -14.99983, 
    -14.99963, -14.99581, 0,
  0, -14.99711, -14.99981, -14.99984, -14.99993, -14.99997, -14.99993, 
    -14.99984, -14.99981, -14.99711, 0,
  0, -14.99999, -14.99988, -14.99989, -14.99984, -14.99983, -14.99984, 
    -14.99989, -14.99988, -14.99999, 0,
  0, -15, -14.99998, -14.99988, -14.99981, -14.99963, -14.99981, -14.99988, 
    -14.99998, -15, 0,
  0, 0, -15, -14.99999, -14.99711, -14.99581, -14.99711, -14.99999, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99998, -14.99215, -14.98863, -14.99215, -14.99998, -15, 0, 0,
  0, -15, -14.99994, -14.99966, -14.99951, -14.99927, -14.99951, -14.99966, 
    -14.99994, -15, 0,
  0, -14.99998, -14.99966, -14.99971, -14.99974, -14.99975, -14.99974, 
    -14.99971, -14.99966, -14.99998, 0,
  0, -14.99215, -14.99951, -14.99974, -14.9999, -14.99996, -14.9999, 
    -14.99974, -14.99951, -14.99215, 0,
  0, -14.98863, -14.99927, -14.99975, -14.99996, -15, -14.99996, -14.99975, 
    -14.99927, -14.98863, 0,
  0, -14.99215, -14.99951, -14.99974, -14.9999, -14.99996, -14.9999, 
    -14.99974, -14.99951, -14.99215, 0,
  0, -14.99998, -14.99966, -14.99971, -14.99974, -14.99975, -14.99974, 
    -14.99971, -14.99966, -14.99998, 0,
  0, -15, -14.99994, -14.99966, -14.99951, -14.99927, -14.99951, -14.99966, 
    -14.99994, -15, 0,
  0, 0, -15, -14.99998, -14.99215, -14.98863, -14.99215, -14.99998, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99994, -14.9883, -14.9831, -14.9883, -14.99994, -15, 0, 0,
  0, -15, -14.99984, -14.99897, -14.99848, -14.99814, -14.99848, -14.99897, 
    -14.99984, -15, 0,
  0, -14.99994, -14.99897, -14.99905, -14.99944, -14.99955, -14.99944, 
    -14.99905, -14.99897, -14.99994, 0,
  0, -14.9883, -14.99848, -14.99944, -14.99985, -14.99995, -14.99985, 
    -14.99944, -14.99848, -14.9883, 0,
  0, -14.9831, -14.99814, -14.99955, -14.99995, -15, -14.99995, -14.99955, 
    -14.99814, -14.9831, 0,
  0, -14.9883, -14.99848, -14.99944, -14.99985, -14.99995, -14.99985, 
    -14.99944, -14.99848, -14.9883, 0,
  0, -14.99994, -14.99897, -14.99905, -14.99944, -14.99955, -14.99944, 
    -14.99905, -14.99897, -14.99994, 0,
  0, -15, -14.99984, -14.99897, -14.99848, -14.99814, -14.99848, -14.99897, 
    -14.99984, -15, 0,
  0, 0, -15, -14.99994, -14.9883, -14.9831, -14.9883, -14.99994, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99989, -14.98517, -14.97866, -14.98517, -14.99989, -15, 0, 0,
  0, -15, -14.99968, -14.99773, -14.9965, -14.99597, -14.9965, -14.99773, 
    -14.99968, -15, 0,
  0, -14.99989, -14.99773, -14.99779, -14.99886, -14.99917, -14.99886, 
    -14.99779, -14.99773, -14.99989, 0,
  0, -14.98517, -14.9965, -14.99886, -14.99977, -14.99993, -14.99977, 
    -14.99886, -14.9965, -14.98517, 0,
  0, -14.97866, -14.99597, -14.99917, -14.99993, -15, -14.99993, -14.99917, 
    -14.99597, -14.97866, 0,
  0, -14.98517, -14.9965, -14.99886, -14.99977, -14.99993, -14.99977, 
    -14.99886, -14.9965, -14.98517, 0,
  0, -14.99989, -14.99773, -14.99779, -14.99886, -14.99917, -14.99886, 
    -14.99779, -14.99773, -14.99989, 0,
  0, -15, -14.99968, -14.99773, -14.9965, -14.99597, -14.9965, -14.99773, 
    -14.99968, -15, 0,
  0, 0, -15, -14.99989, -14.98517, -14.97866, -14.98517, -14.99989, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99983, -14.98267, -14.97501, -14.98267, -14.99983, -15, 0, 0,
  0, -15, -14.99948, -14.99582, -14.99374, -14.99291, -14.99374, -14.99582, 
    -14.99948, -15, 0,
  0, -14.99983, -14.99582, -14.99604, -14.99806, -14.99864, -14.99806, 
    -14.99604, -14.99582, -14.99983, 0,
  0, -14.98267, -14.99374, -14.99806, -14.99965, -14.9999, -14.99965, 
    -14.99806, -14.99374, -14.98267, 0,
  0, -14.97501, -14.99291, -14.99864, -14.9999, -15, -14.9999, -14.99864, 
    -14.99291, -14.97501, 0,
  0, -14.98267, -14.99374, -14.99806, -14.99965, -14.9999, -14.99965, 
    -14.99806, -14.99374, -14.98267, 0,
  0, -14.99983, -14.99582, -14.99604, -14.99806, -14.99864, -14.99806, 
    -14.99604, -14.99582, -14.99983, 0,
  0, -15, -14.99948, -14.99582, -14.99374, -14.99291, -14.99374, -14.99582, 
    -14.99948, -15, 0,
  0, 0, -15, -14.99983, -14.98267, -14.97501, -14.98267, -14.99983, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99971, -14.98061, -14.97207, -14.98061, -14.99971, -15, 0, 0,
  0, -15, -14.99907, -14.99147, -14.99024, -14.98911, -14.99024, -14.99147, 
    -14.99907, -15, 0,
  0, -14.99971, -14.99147, -14.99387, -14.99707, -14.99798, -14.99707, 
    -14.99387, -14.99147, -14.99971, 0,
  0, -14.98061, -14.99024, -14.99707, -14.99949, -14.99984, -14.99949, 
    -14.99707, -14.99024, -14.98061, 0,
  0, -14.97207, -14.98911, -14.99798, -14.99984, -14.99999, -14.99984, 
    -14.99798, -14.98911, -14.97207, 0,
  0, -14.98061, -14.99024, -14.99707, -14.99949, -14.99984, -14.99949, 
    -14.99707, -14.99024, -14.98061, 0,
  0, -14.99971, -14.99147, -14.99387, -14.99707, -14.99798, -14.99707, 
    -14.99387, -14.99147, -14.99971, 0,
  0, -15, -14.99907, -14.99147, -14.99024, -14.98911, -14.99024, -14.99147, 
    -14.99907, -15, 0,
  0, 0, -15, -14.99971, -14.98061, -14.97207, -14.98061, -14.99971, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99934, -14.97885, -14.96959, -14.97885, -14.99934, -15, 0, 0,
  0, -15, -14.99753, -14.97532, -14.98331, -14.9827, -14.98331, -14.97532, 
    -14.99753, -15, 0,
  0, -14.99934, -14.97532, -14.98981, -14.99514, -14.99654, -14.99514, 
    -14.98981, -14.97532, -14.99934, 0,
  0, -14.97885, -14.98331, -14.99514, -14.99881, -14.99937, -14.99881, 
    -14.99514, -14.98331, -14.97885, 0,
  0, -14.96959, -14.9827, -14.99654, -14.99937, -14.99962, -14.99937, 
    -14.99654, -14.9827, -14.96959, 0,
  0, -14.97885, -14.98331, -14.99514, -14.99881, -14.99937, -14.99881, 
    -14.99514, -14.98331, -14.97885, 0,
  0, -14.99934, -14.97532, -14.98981, -14.99514, -14.99654, -14.99514, 
    -14.98981, -14.97532, -14.99934, 0,
  0, -15, -14.99753, -14.97532, -14.98331, -14.9827, -14.98331, -14.97532, 
    -14.99753, -15, 0,
  0, 0, -15, -14.99934, -14.97885, -14.96959, -14.97885, -14.99934, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.9987, -14.97719, -14.96737, -14.97719, -14.9987, -15, 0, 0,
  0, -15, -14.99424, -14.91986, -14.95236, -14.95567, -14.95236, -14.91986, 
    -14.99424, -15, 0,
  0, -14.9987, -14.91986, -14.96781, -14.98072, -14.98386, -14.98072, 
    -14.96781, -14.91986, -14.9987, 0,
  0, -14.97719, -14.95236, -14.98072, -14.98891, -14.99047, -14.98891, 
    -14.98072, -14.95236, -14.97719, 0,
  0, -14.96737, -14.95567, -14.98386, -14.99047, -14.99153, -14.99047, 
    -14.98386, -14.95567, -14.96737, 0,
  0, -14.97719, -14.95236, -14.98072, -14.98891, -14.99047, -14.98891, 
    -14.98072, -14.95236, -14.97719, 0,
  0, -14.9987, -14.91986, -14.96781, -14.98072, -14.98386, -14.98072, 
    -14.96781, -14.91986, -14.9987, 0,
  0, -15, -14.99424, -14.91986, -14.95236, -14.95567, -14.95236, -14.91986, 
    -14.99424, -15, 0,
  0, 0, -15, -14.9987, -14.97719, -14.96737, -14.97719, -14.9987, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99877, -14.97582, -14.96538, -14.97582, -14.99877, -15, 0, 0,
  0, -15, -14.99318, -14.7823, -14.81684, -14.8234, -14.81684, -14.7823, 
    -14.99318, -15, 0,
  0, -14.99877, -14.7823, -14.8404, -14.86465, -14.87114, -14.86465, 
    -14.8404, -14.7823, -14.99877, 0,
  0, -14.97582, -14.81684, -14.86465, -14.88219, -14.88636, -14.88219, 
    -14.86465, -14.81684, -14.97582, 0,
  0, -14.96538, -14.8234, -14.87114, -14.88636, -14.8898, -14.88636, 
    -14.87114, -14.8234, -14.96538, 0,
  0, -14.97582, -14.81684, -14.86465, -14.88219, -14.88636, -14.88219, 
    -14.86465, -14.81684, -14.97582, 0,
  0, -14.99877, -14.7823, -14.8404, -14.86465, -14.87114, -14.86465, 
    -14.8404, -14.7823, -14.99877, 0,
  0, -15, -14.99318, -14.7823, -14.81684, -14.8234, -14.81684, -14.7823, 
    -14.99318, -15, 0,
  0, 0, -15, -14.99877, -14.97582, -14.96538, -14.97582, -14.99877, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -14.97585, -14.96517, -14.97585, -15, -15, -15, -15,
  -15, -15, -15, -14.65447, -14.61903, -14.6074, -14.61903, -14.65447, -15, 
    -15, -15,
  -15, -15, -14.65447, -14.60733, -14.58711, -14.58027, -14.58711, -14.60733, 
    -14.65447, -15, -15,
  -15, -14.97585, -14.61903, -14.58711, -14.56597, -14.55814, -14.56597, 
    -14.58711, -14.61903, -14.97585, -15,
  -15, -14.96517, -14.6074, -14.58027, -14.55814, -14.55001, -14.55814, 
    -14.58027, -14.6074, -14.96517, -15,
  -15, -14.97585, -14.61903, -14.58711, -14.56597, -14.55814, -14.56597, 
    -14.58711, -14.61903, -14.97585, -15,
  -15, -15, -14.65447, -14.60733, -14.58711, -14.58027, -14.58711, -14.60733, 
    -14.65447, -15, -15,
  -15, -15, -15, -14.65447, -14.61903, -14.6074, -14.61903, -14.65447, -15, 
    -15, -15,
  -15, -15, -15, -15, -14.97585, -14.96517, -14.97585, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99999, -14.99692, -14.99559, -14.99692, -14.99999, -15, 0, 0,
  0, -15, -14.99998, -14.99985, -14.99979, -14.99961, -14.99979, -14.99985, 
    -14.99998, -15, 0,
  0, -14.99999, -14.99985, -14.99986, -14.9998, -14.99979, -14.9998, 
    -14.99986, -14.99985, -14.99999, 0,
  0, -14.99692, -14.99979, -14.9998, -14.99991, -14.99996, -14.99991, 
    -14.9998, -14.99979, -14.99692, 0,
  0, -14.99559, -14.99961, -14.99979, -14.99996, -15, -14.99996, -14.99979, 
    -14.99961, -14.99559, 0,
  0, -14.99692, -14.99979, -14.9998, -14.99991, -14.99996, -14.99991, 
    -14.9998, -14.99979, -14.99692, 0,
  0, -14.99999, -14.99985, -14.99986, -14.9998, -14.99979, -14.9998, 
    -14.99986, -14.99985, -14.99999, 0,
  0, -15, -14.99998, -14.99985, -14.99979, -14.99961, -14.99979, -14.99985, 
    -14.99998, -15, 0,
  0, 0, -15, -14.99999, -14.99692, -14.99559, -14.99692, -14.99999, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99997, -14.99165, -14.98803, -14.99165, -14.99997, -15, 0, 0,
  0, -15, -14.99994, -14.99958, -14.99945, -14.99921, -14.99945, -14.99958, 
    -14.99994, -15, 0,
  0, -14.99997, -14.99958, -14.99963, -14.99968, -14.9997, -14.99968, 
    -14.99963, -14.99958, -14.99997, 0,
  0, -14.99165, -14.99945, -14.99968, -14.99988, -14.99995, -14.99988, 
    -14.99968, -14.99945, -14.99165, 0,
  0, -14.98803, -14.99921, -14.9997, -14.99995, -15, -14.99995, -14.9997, 
    -14.99921, -14.98803, 0,
  0, -14.99165, -14.99945, -14.99968, -14.99988, -14.99995, -14.99988, 
    -14.99968, -14.99945, -14.99165, 0,
  0, -14.99997, -14.99958, -14.99963, -14.99968, -14.9997, -14.99968, 
    -14.99963, -14.99958, -14.99997, 0,
  0, -15, -14.99994, -14.99958, -14.99945, -14.99921, -14.99945, -14.99958, 
    -14.99994, -15, 0,
  0, 0, -15, -14.99997, -14.99165, -14.98803, -14.99165, -14.99997, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99993, -14.98755, -14.98222, -14.98755, -14.99993, -15, 0, 0,
  0, -15, -14.99983, -14.99877, -14.99829, -14.99796, -14.99829, -14.99877, 
    -14.99983, -15, 0,
  0, -14.99993, -14.99877, -14.99882, -14.99931, -14.99945, -14.99931, 
    -14.99882, -14.99877, -14.99993, 0,
  0, -14.98755, -14.99829, -14.99931, -14.99982, -14.99993, -14.99982, 
    -14.99931, -14.99829, -14.98755, 0,
  0, -14.98222, -14.99796, -14.99945, -14.99993, -15, -14.99993, -14.99945, 
    -14.99796, -14.98222, 0,
  0, -14.98755, -14.99829, -14.99931, -14.99982, -14.99993, -14.99982, 
    -14.99931, -14.99829, -14.98755, 0,
  0, -14.99993, -14.99877, -14.99882, -14.99931, -14.99945, -14.99931, 
    -14.99882, -14.99877, -14.99993, 0,
  0, -15, -14.99983, -14.99877, -14.99829, -14.99796, -14.99829, -14.99877, 
    -14.99983, -15, 0,
  0, 0, -15, -14.99993, -14.98755, -14.98222, -14.98755, -14.99993, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99987, -14.98425, -14.97755, -14.98425, -14.99987, -15, 0, 0,
  0, -15, -14.99967, -14.99727, -14.99607, -14.99555, -14.99607, -14.99727, 
    -14.99967, -15, 0,
  0, -14.99987, -14.99727, -14.99726, -14.9986, -14.99898, -14.9986, 
    -14.99726, -14.99727, -14.99987, 0,
  0, -14.98425, -14.99607, -14.9986, -14.99971, -14.99991, -14.99971, 
    -14.9986, -14.99607, -14.98425, 0,
  0, -14.97755, -14.99555, -14.99898, -14.99991, -15, -14.99991, -14.99898, 
    -14.99555, -14.97755, 0,
  0, -14.98425, -14.99607, -14.9986, -14.99971, -14.99991, -14.99971, 
    -14.9986, -14.99607, -14.98425, 0,
  0, -14.99987, -14.99727, -14.99726, -14.9986, -14.99898, -14.9986, 
    -14.99726, -14.99727, -14.99987, 0,
  0, -15, -14.99967, -14.99727, -14.99607, -14.99555, -14.99607, -14.99727, 
    -14.99967, -15, 0,
  0, 0, -15, -14.99987, -14.98425, -14.97755, -14.98425, -14.99987, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.9998, -14.98161, -14.97374, -14.98161, -14.9998, -15, 0, 0,
  0, -15, -14.99944, -14.9948, -14.99298, -14.99216, -14.99298, -14.9948, 
    -14.99944, -15, 0,
  0, -14.9998, -14.9948, -14.99507, -14.9976, -14.99832, -14.9976, -14.99507, 
    -14.9948, -14.9998, 0,
  0, -14.98161, -14.99298, -14.9976, -14.99956, -14.99987, -14.99956, 
    -14.9976, -14.99298, -14.98161, 0,
  0, -14.97374, -14.99216, -14.99832, -14.99987, -15, -14.99987, -14.99832, 
    -14.99216, -14.97374, 0,
  0, -14.98161, -14.99298, -14.9976, -14.99956, -14.99987, -14.99956, 
    -14.9976, -14.99298, -14.98161, 0,
  0, -14.9998, -14.9948, -14.99507, -14.9976, -14.99832, -14.9976, -14.99507, 
    -14.9948, -14.9998, 0,
  0, -15, -14.99944, -14.9948, -14.99298, -14.99216, -14.99298, -14.9948, 
    -14.99944, -15, 0,
  0, 0, -15, -14.9998, -14.98161, -14.97374, -14.98161, -14.9998, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99963, -14.97944, -14.97066, -14.97944, -14.99963, -15, 0, 0,
  0, -15, -14.99891, -14.98845, -14.98887, -14.98784, -14.98887, -14.98845, 
    -14.99891, -15, 0,
  0, -14.99963, -14.98845, -14.99231, -14.99634, -14.99748, -14.99634, 
    -14.99231, -14.98845, -14.99963, 0,
  0, -14.97944, -14.98887, -14.99634, -14.99934, -14.9998, -14.99934, 
    -14.99634, -14.98887, -14.97944, 0,
  0, -14.97066, -14.98784, -14.99748, -14.9998, -14.99998, -14.9998, 
    -14.99748, -14.98784, -14.97066, 0,
  0, -14.97944, -14.98887, -14.99634, -14.99934, -14.9998, -14.99934, 
    -14.99634, -14.98887, -14.97944, 0,
  0, -14.99963, -14.98845, -14.99231, -14.99634, -14.99748, -14.99634, 
    -14.99231, -14.98845, -14.99963, 0,
  0, -15, -14.99891, -14.98845, -14.98887, -14.98784, -14.98887, -14.98845, 
    -14.99891, -15, 0,
  0, 0, -15, -14.99963, -14.97944, -14.97066, -14.97944, -14.99963, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99912, -14.97757, -14.96805, -14.97757, -14.99912, -15, 0, 0,
  0, -15, -14.99707, -14.9655, -14.9795, -14.97952, -14.9795, -14.9655, 
    -14.99707, -15, 0,
  0, -14.99912, -14.9655, -14.98655, -14.99356, -14.99538, -14.99356, 
    -14.98655, -14.9655, -14.99912, 0,
  0, -14.97757, -14.9795, -14.99356, -14.99828, -14.99901, -14.99828, 
    -14.99356, -14.9795, -14.97757, 0,
  0, -14.96805, -14.97952, -14.99538, -14.99901, -14.99936, -14.99901, 
    -14.99538, -14.97952, -14.96805, 0,
  0, -14.97757, -14.9795, -14.99356, -14.99828, -14.99901, -14.99828, 
    -14.99356, -14.9795, -14.97757, 0,
  0, -14.99912, -14.9655, -14.98655, -14.99356, -14.99538, -14.99356, 
    -14.98655, -14.9655, -14.99912, 0,
  0, -15, -14.99707, -14.9655, -14.9795, -14.97952, -14.9795, -14.9655, 
    -14.99707, -15, 0,
  0, 0, -15, -14.99912, -14.97757, -14.96805, -14.97757, -14.99912, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99838, -14.97576, -14.96566, -14.97576, -14.99838, -15, 0, 0,
  0, -15, -14.99386, -14.89564, -14.93822, -14.94335, -14.93822, -14.89564, 
    -14.99386, -15, 0,
  0, -14.99838, -14.89564, -14.95624, -14.97326, -14.97741, -14.97326, 
    -14.95624, -14.89564, -14.99838, 0,
  0, -14.97576, -14.93822, -14.97326, -14.98408, -14.9862, -14.98408, 
    -14.97326, -14.93822, -14.97576, 0,
  0, -14.96566, -14.94335, -14.97741, -14.9862, -14.98767, -14.9862, 
    -14.97741, -14.94335, -14.96566, 0,
  0, -14.97576, -14.93822, -14.97326, -14.98408, -14.9862, -14.98408, 
    -14.97326, -14.93822, -14.97576, 0,
  0, -14.99838, -14.89564, -14.95624, -14.97326, -14.97741, -14.97326, 
    -14.95624, -14.89564, -14.99838, 0,
  0, -15, -14.99386, -14.89564, -14.93822, -14.94335, -14.93822, -14.89564, 
    -14.99386, -15, 0,
  0, 0, -15, -14.99838, -14.97576, -14.96566, -14.97576, -14.99838, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99861, -14.97436, -14.96361, -14.97436, -14.99861, -15, 0, 0,
  0, -15, -14.99375, -14.74352, -14.78144, -14.78908, -14.78144, -14.74352, 
    -14.99375, -15, 0,
  0, -14.99861, -14.74352, -14.80617, -14.8346, -14.84231, -14.8346, 
    -14.80617, -14.74352, -14.99861, 0,
  0, -14.97436, -14.78144, -14.8346, -14.85548, -14.86047, -14.85548, 
    -14.8346, -14.78144, -14.97436, 0,
  0, -14.96361, -14.78908, -14.84231, -14.86047, -14.86457, -14.86047, 
    -14.84231, -14.78908, -14.96361, 0,
  0, -14.97436, -14.78144, -14.8346, -14.85548, -14.86047, -14.85548, 
    -14.8346, -14.78144, -14.97436, 0,
  0, -14.99861, -14.74352, -14.80617, -14.8346, -14.84231, -14.8346, 
    -14.80617, -14.74352, -14.99861, 0,
  0, -15, -14.99375, -14.74352, -14.78144, -14.78908, -14.78144, -14.74352, 
    -14.99375, -15, 0,
  0, 0, -15, -14.99861, -14.97436, -14.96361, -14.97436, -14.99861, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -14.97447, -14.96348, -14.97447, -15, -15, -15, -15,
  -15, -15, -15, -14.61556, -14.58351, -14.57296, -14.58351, -14.61556, -15, 
    -15, -15,
  -15, -15, -14.61556, -14.57315, -14.55722, -14.55162, -14.55722, -14.57315, 
    -14.61556, -15, -15,
  -15, -14.97447, -14.58351, -14.55722, -14.53937, -14.53231, -14.53937, 
    -14.55722, -14.58351, -14.97447, -15,
  -15, -14.96348, -14.57296, -14.55162, -14.53231, -14.52479, -14.53231, 
    -14.55162, -14.57296, -14.96348, -15,
  -15, -14.97447, -14.58351, -14.55722, -14.53937, -14.53231, -14.53937, 
    -14.55722, -14.58351, -14.97447, -15,
  -15, -15, -14.61556, -14.57315, -14.55722, -14.55162, -14.55722, -14.57315, 
    -14.61556, -15, -15,
  -15, -15, -15, -14.61556, -14.58351, -14.57296, -14.58351, -14.61556, -15, 
    -15, -15,
  -15, -15, -15, -15, -14.97447, -14.96348, -14.97447, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99999, -14.99677, -14.99539, -14.99677, -14.99999, -15, 0, 0,
  0, -15, -14.99997, -14.99981, -14.99976, -14.99959, -14.99976, -14.99981, 
    -14.99997, -15, 0,
  0, -14.99999, -14.99981, -14.99984, -14.99977, -14.99975, -14.99977, 
    -14.99984, -14.99981, -14.99999, 0,
  0, -14.99677, -14.99976, -14.99977, -14.99989, -14.99995, -14.99989, 
    -14.99977, -14.99976, -14.99677, 0,
  0, -14.99539, -14.99959, -14.99975, -14.99995, -15, -14.99995, -14.99975, 
    -14.99959, -14.99539, 0,
  0, -14.99677, -14.99976, -14.99977, -14.99989, -14.99995, -14.99989, 
    -14.99977, -14.99976, -14.99677, 0,
  0, -14.99999, -14.99981, -14.99984, -14.99977, -14.99975, -14.99977, 
    -14.99984, -14.99981, -14.99999, 0,
  0, -15, -14.99997, -14.99981, -14.99976, -14.99959, -14.99976, -14.99981, 
    -14.99997, -15, 0,
  0, 0, -15, -14.99999, -14.99677, -14.99539, -14.99677, -14.99999, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99997, -14.99123, -14.98748, -14.99123, -14.99997, -15, 0, 0,
  0, -15, -14.99993, -14.9995, -14.99938, -14.99915, -14.99938, -14.9995, 
    -14.99993, -15, 0,
  0, -14.99997, -14.9995, -14.99956, -14.99962, -14.99965, -14.99962, 
    -14.99956, -14.9995, -14.99997, 0,
  0, -14.99123, -14.99938, -14.99962, -14.99985, -14.99994, -14.99985, 
    -14.99962, -14.99938, -14.99123, 0,
  0, -14.98748, -14.99915, -14.99965, -14.99994, -15, -14.99994, -14.99965, 
    -14.99915, -14.98748, 0,
  0, -14.99123, -14.99938, -14.99962, -14.99985, -14.99994, -14.99985, 
    -14.99962, -14.99938, -14.99123, 0,
  0, -14.99997, -14.9995, -14.99956, -14.99962, -14.99965, -14.99962, 
    -14.99956, -14.9995, -14.99997, 0,
  0, -15, -14.99993, -14.9995, -14.99938, -14.99915, -14.99938, -14.9995, 
    -14.99993, -15, 0,
  0, 0, -15, -14.99997, -14.99123, -14.98748, -14.99123, -14.99997, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99993, -14.98694, -14.9814, -14.98694, -14.99993, -15, 0, 0,
  0, -15, -14.99982, -14.99855, -14.9981, -14.99778, -14.9981, -14.99855, 
    -14.99982, -15, 0,
  0, -14.99993, -14.99855, -14.99859, -14.99918, -14.99935, -14.99918, 
    -14.99859, -14.99855, -14.99993, 0,
  0, -14.98694, -14.9981, -14.99918, -14.99978, -14.99992, -14.99978, 
    -14.99918, -14.9981, -14.98694, 0,
  0, -14.9814, -14.99778, -14.99935, -14.99992, -15, -14.99992, -14.99935, 
    -14.99778, -14.9814, 0,
  0, -14.98694, -14.9981, -14.99918, -14.99978, -14.99992, -14.99978, 
    -14.99918, -14.9981, -14.98694, 0,
  0, -14.99993, -14.99855, -14.99859, -14.99918, -14.99935, -14.99918, 
    -14.99859, -14.99855, -14.99993, 0,
  0, -15, -14.99982, -14.99855, -14.9981, -14.99778, -14.9981, -14.99855, 
    -14.99982, -15, 0,
  0, 0, -15, -14.99993, -14.98694, -14.9814, -14.98694, -14.99993, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99986, -14.98348, -14.97652, -14.98348, -14.99986, -15, 0, 0,
  0, -15, -14.99965, -14.99679, -14.99565, -14.99513, -14.99565, -14.99679, 
    -14.99965, -15, 0,
  0, -14.99986, -14.99679, -14.99672, -14.99833, -14.99879, -14.99833, 
    -14.99672, -14.99679, -14.99986, 0,
  0, -14.98348, -14.99565, -14.99833, -14.99965, -14.99989, -14.99965, 
    -14.99833, -14.99565, -14.98348, 0,
  0, -14.97652, -14.99513, -14.99879, -14.99989, -15, -14.99989, -14.99879, 
    -14.99513, -14.97652, 0,
  0, -14.98348, -14.99565, -14.99833, -14.99965, -14.99989, -14.99965, 
    -14.99833, -14.99565, -14.98348, 0,
  0, -14.99986, -14.99679, -14.99672, -14.99833, -14.99879, -14.99833, 
    -14.99672, -14.99679, -14.99986, 0,
  0, -15, -14.99965, -14.99679, -14.99565, -14.99513, -14.99565, -14.99679, 
    -14.99965, -15, 0,
  0, 0, -15, -14.99986, -14.98348, -14.97652, -14.98348, -14.99986, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99977, -14.98072, -14.97254, -14.98072, -14.99977, -15, 0, 0,
  0, -15, -14.99939, -14.99364, -14.99221, -14.9914, -14.99221, -14.99364, 
    -14.99939, -15, 0,
  0, -14.99977, -14.99364, -14.99411, -14.99714, -14.998, -14.99714, 
    -14.99411, -14.99364, -14.99977, 0,
  0, -14.98072, -14.99221, -14.99714, -14.99946, -14.99984, -14.99946, 
    -14.99714, -14.99221, -14.98072, 0,
  0, -14.97254, -14.9914, -14.998, -14.99984, -15, -14.99984, -14.998, 
    -14.9914, -14.97254, 0,
  0, -14.98072, -14.99221, -14.99714, -14.99946, -14.99984, -14.99946, 
    -14.99714, -14.99221, -14.98072, 0,
  0, -14.99977, -14.99364, -14.99411, -14.99714, -14.998, -14.99714, 
    -14.99411, -14.99364, -14.99977, 0,
  0, -15, -14.99939, -14.99364, -14.99221, -14.9914, -14.99221, -14.99364, 
    -14.99939, -15, 0,
  0, 0, -15, -14.99977, -14.98072, -14.97254, -14.98072, -14.99977, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99954, -14.97844, -14.96933, -14.97844, -14.99954, -15, 0, 0,
  0, -15, -14.99873, -14.98483, -14.9874, -14.9865, -14.9874, -14.98483, 
    -14.99873, -15, 0,
  0, -14.99954, -14.98483, -14.99071, -14.9956, -14.99697, -14.9956, 
    -14.99071, -14.98483, -14.99954, 0,
  0, -14.97844, -14.9874, -14.9956, -14.99919, -14.99974, -14.99919, 
    -14.9956, -14.9874, -14.97844, 0,
  0, -14.96933, -14.9865, -14.99697, -14.99974, -14.99996, -14.99974, 
    -14.99697, -14.9865, -14.96933, 0,
  0, -14.97844, -14.9874, -14.9956, -14.99919, -14.99974, -14.99919, 
    -14.9956, -14.9874, -14.97844, 0,
  0, -14.99954, -14.98483, -14.99071, -14.9956, -14.99697, -14.9956, 
    -14.99071, -14.98483, -14.99954, 0,
  0, -15, -14.99873, -14.98483, -14.9874, -14.9865, -14.9874, -14.98483, 
    -14.99873, -15, 0,
  0, 0, -15, -14.99954, -14.97844, -14.96933, -14.97844, -14.99954, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99889, -14.97646, -14.96659, -14.97646, -14.99889, -15, 0, 0,
  0, -15, -14.99665, -14.95452, -14.97513, -14.97589, -14.97513, -14.95452, 
    -14.99665, -15, 0,
  0, -14.99889, -14.95452, -14.98294, -14.99178, -14.99404, -14.99178, 
    -14.98294, -14.95452, -14.99889, 0,
  0, -14.97646, -14.97513, -14.99178, -14.99762, -14.99855, -14.99762, 
    -14.99178, -14.97513, -14.97646, 0,
  0, -14.96659, -14.97589, -14.99404, -14.99855, -14.99901, -14.99855, 
    -14.99404, -14.97589, -14.96659, 0,
  0, -14.97646, -14.97513, -14.99178, -14.99762, -14.99855, -14.99762, 
    -14.99178, -14.97513, -14.97646, 0,
  0, -14.99889, -14.95452, -14.98294, -14.99178, -14.99404, -14.99178, 
    -14.98294, -14.95452, -14.99889, 0,
  0, -15, -14.99665, -14.95452, -14.97513, -14.97589, -14.97513, -14.95452, 
    -14.99665, -15, 0,
  0, 0, -15, -14.99889, -14.97646, -14.96659, -14.97646, -14.99889, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99808, -14.97452, -14.96405, -14.97452, -14.99808, -15, 0, 0,
  0, -15, -14.99359, -14.87141, -14.92318, -14.93012, -14.92318, -14.87141, 
    -14.99359, -15, 0,
  0, -14.99808, -14.87141, -14.94376, -14.96501, -14.97022, -14.96501, 
    -14.94376, -14.87141, -14.99808, 0,
  0, -14.97452, -14.92318, -14.96501, -14.9786, -14.98132, -14.9786, 
    -14.96501, -14.92318, -14.97452, 0,
  0, -14.96405, -14.93012, -14.97022, -14.98132, -14.98325, -14.98132, 
    -14.97022, -14.93012, -14.96405, 0,
  0, -14.97452, -14.92318, -14.96501, -14.9786, -14.98132, -14.9786, 
    -14.96501, -14.92318, -14.97452, 0,
  0, -14.99808, -14.87141, -14.94376, -14.96501, -14.97022, -14.96501, 
    -14.94376, -14.87141, -14.99808, 0,
  0, -15, -14.99359, -14.87141, -14.92318, -14.93012, -14.92318, -14.87141, 
    -14.99359, -15, 0,
  0, 0, -15, -14.99808, -14.97452, -14.96405, -14.97452, -14.99808, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99848, -14.97309, -14.96194, -14.97309, -14.99848, -15, 0, 0,
  0, -15, -14.99418, -14.70796, -14.74823, -14.7567, -14.74823, -14.70796, 
    -14.99418, -15, 0,
  0, -14.99848, -14.70796, -14.77366, -14.80581, -14.81461, -14.80581, 
    -14.77366, -14.70796, -14.99848, 0,
  0, -14.97309, -14.74823, -14.80581, -14.82972, -14.83545, -14.82972, 
    -14.80581, -14.74823, -14.97309, 0,
  0, -14.96194, -14.7567, -14.81461, -14.83545, -14.84016, -14.83545, 
    -14.81461, -14.7567, -14.96194, 0,
  0, -14.97309, -14.74823, -14.80581, -14.82972, -14.83545, -14.82972, 
    -14.80581, -14.74823, -14.97309, 0,
  0, -14.99848, -14.70796, -14.77366, -14.80581, -14.81461, -14.80581, 
    -14.77366, -14.70796, -14.99848, 0,
  0, -15, -14.99418, -14.70796, -14.74823, -14.7567, -14.74823, -14.70796, 
    -14.99418, -15, 0,
  0, 0, -15, -14.99848, -14.97309, -14.96194, -14.97309, -14.99848, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -14.97327, -14.96187, -14.97327, -15, -15, -15, -15,
  -15, -15, -15, -14.57988, -14.55017, -14.54046, -14.55017, -14.57988, -15, 
    -15, -15,
  -15, -15, -14.57988, -14.5407, -14.52857, -14.52409, -14.52857, -14.5407, 
    -14.57988, -15, -15,
  -15, -14.97327, -14.55017, -14.52857, -14.51372, -14.50735, -14.51372, 
    -14.52857, -14.55017, -14.97327, -15,
  -15, -14.96187, -14.54046, -14.52409, -14.50735, -14.50039, -14.50735, 
    -14.52409, -14.54046, -14.96187, -15,
  -15, -14.97327, -14.55017, -14.52857, -14.51372, -14.50735, -14.51372, 
    -14.52857, -14.55017, -14.97327, -15,
  -15, -15, -14.57988, -14.5407, -14.52857, -14.52409, -14.52857, -14.5407, 
    -14.57988, -15, -15,
  -15, -15, -15, -14.57988, -14.55017, -14.54046, -14.55017, -14.57988, -15, 
    -15, -15,
  -15, -15, -15, -15, -14.97327, -14.96187, -14.97327, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99999, -14.99662, -14.99519, -14.99662, -14.99999, -15, 0, 0,
  0, -15, -14.99997, -14.99978, -14.99974, -14.99957, -14.99974, -14.99978, 
    -14.99997, -15, 0,
  0, -14.99999, -14.99978, -14.99981, -14.99973, -14.99972, -14.99973, 
    -14.99981, -14.99978, -14.99999, 0,
  0, -14.99662, -14.99974, -14.99973, -14.99987, -14.99995, -14.99987, 
    -14.99973, -14.99974, -14.99662, 0,
  0, -14.99519, -14.99957, -14.99972, -14.99995, -15, -14.99995, -14.99972, 
    -14.99957, -14.99519, 0,
  0, -14.99662, -14.99974, -14.99973, -14.99987, -14.99995, -14.99987, 
    -14.99973, -14.99974, -14.99662, 0,
  0, -14.99999, -14.99978, -14.99981, -14.99973, -14.99972, -14.99973, 
    -14.99981, -14.99978, -14.99999, 0,
  0, -15, -14.99997, -14.99978, -14.99974, -14.99957, -14.99974, -14.99978, 
    -14.99997, -15, 0,
  0, 0, -15, -14.99999, -14.99662, -14.99519, -14.99662, -14.99999, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99997, -14.99082, -14.98692, -14.99082, -14.99997, -15, 0, 0,
  0, -15, -14.99993, -14.99942, -14.99932, -14.99909, -14.99932, -14.99942, 
    -14.99993, -15, 0,
  0, -14.99997, -14.99942, -14.99948, -14.99956, -14.99959, -14.99956, 
    -14.99948, -14.99942, -14.99997, 0,
  0, -14.99082, -14.99932, -14.99956, -14.99983, -14.99993, -14.99983, 
    -14.99956, -14.99932, -14.99082, 0,
  0, -14.98692, -14.99909, -14.99959, -14.99993, -15, -14.99993, -14.99959, 
    -14.99909, -14.98692, 0,
  0, -14.99082, -14.99932, -14.99956, -14.99983, -14.99993, -14.99983, 
    -14.99956, -14.99932, -14.99082, 0,
  0, -14.99997, -14.99942, -14.99948, -14.99956, -14.99959, -14.99956, 
    -14.99948, -14.99942, -14.99997, 0,
  0, -15, -14.99993, -14.99942, -14.99932, -14.99909, -14.99932, -14.99942, 
    -14.99993, -15, 0,
  0, 0, -15, -14.99997, -14.99082, -14.98692, -14.99082, -14.99997, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99992, -14.98632, -14.98057, -14.98632, -14.99992, -15, 0, 0,
  0, -15, -14.99982, -14.99833, -14.99791, -14.99759, -14.99791, -14.99833, 
    -14.99982, -15, 0,
  0, -14.99992, -14.99833, -14.99836, -14.99905, -14.99925, -14.99905, 
    -14.99836, -14.99833, -14.99992, 0,
  0, -14.98632, -14.99791, -14.99905, -14.99974, -14.9999, -14.99974, 
    -14.99905, -14.99791, -14.98632, 0,
  0, -14.98057, -14.99759, -14.99925, -14.9999, -15, -14.9999, -14.99925, 
    -14.99759, -14.98057, 0,
  0, -14.98632, -14.99791, -14.99905, -14.99974, -14.9999, -14.99974, 
    -14.99905, -14.99791, -14.98632, 0,
  0, -14.99992, -14.99833, -14.99836, -14.99905, -14.99925, -14.99905, 
    -14.99836, -14.99833, -14.99992, 0,
  0, -15, -14.99982, -14.99833, -14.99791, -14.99759, -14.99791, -14.99833, 
    -14.99982, -15, 0,
  0, 0, -15, -14.99992, -14.98632, -14.98057, -14.98632, -14.99992, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99985, -14.98271, -14.97548, -14.98271, -14.99985, -15, 0, 0,
  0, -15, -14.99964, -14.99628, -14.99522, -14.99471, -14.99522, -14.99628, 
    -14.99964, -15, 0,
  0, -14.99985, -14.99628, -14.99618, -14.99806, -14.99861, -14.99806, 
    -14.99618, -14.99628, -14.99985, 0,
  0, -14.98271, -14.99522, -14.99806, -14.99959, -14.99987, -14.99959, 
    -14.99806, -14.99522, -14.98271, 0,
  0, -14.97548, -14.99471, -14.99861, -14.99987, -15, -14.99987, -14.99861, 
    -14.99471, -14.97548, 0,
  0, -14.98271, -14.99522, -14.99806, -14.99959, -14.99987, -14.99959, 
    -14.99806, -14.99522, -14.98271, 0,
  0, -14.99985, -14.99628, -14.99618, -14.99806, -14.99861, -14.99806, 
    -14.99618, -14.99628, -14.99985, 0,
  0, -15, -14.99964, -14.99628, -14.99522, -14.99471, -14.99522, -14.99628, 
    -14.99964, -15, 0,
  0, 0, -15, -14.99985, -14.98271, -14.97548, -14.98271, -14.99985, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99973, -14.97983, -14.97134, -14.97983, -14.99973, -15, 0, 0,
  0, -15, -14.99934, -14.99233, -14.99142, -14.99064, -14.99142, -14.99233, 
    -14.99934, -15, 0,
  0, -14.99973, -14.99233, -14.99314, -14.99667, -14.99769, -14.99667, 
    -14.99314, -14.99233, -14.99973, 0,
  0, -14.97983, -14.99142, -14.99667, -14.99937, -14.99981, -14.99937, 
    -14.99667, -14.99142, -14.97983, 0,
  0, -14.97134, -14.99064, -14.99769, -14.99981, -15, -14.99981, -14.99769, 
    -14.99064, -14.97134, 0,
  0, -14.97983, -14.99142, -14.99667, -14.99937, -14.99981, -14.99937, 
    -14.99667, -14.99142, -14.97983, 0,
  0, -14.99973, -14.99233, -14.99314, -14.99667, -14.99769, -14.99667, 
    -14.99314, -14.99233, -14.99973, 0,
  0, -15, -14.99934, -14.99233, -14.99142, -14.99064, -14.99142, -14.99233, 
    -14.99934, -15, 0,
  0, 0, -15, -14.99973, -14.97983, -14.97134, -14.97983, -14.99973, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.9994, -14.97744, -14.96799, -14.97744, -14.9994, -15, 0, 0,
  0, -15, -14.99846, -14.98064, -14.98581, -14.98509, -14.98581, -14.98064, 
    -14.99846, -15, 0,
  0, -14.9994, -14.98064, -14.98906, -14.99483, -14.99644, -14.99483, 
    -14.98906, -14.98064, -14.9994, 0,
  0, -14.97744, -14.98581, -14.99483, -14.99903, -14.99967, -14.99903, 
    -14.99483, -14.98581, -14.97744, 0,
  0, -14.96799, -14.98509, -14.99644, -14.99967, -14.99994, -14.99967, 
    -14.99644, -14.98509, -14.96799, 0,
  0, -14.97744, -14.98581, -14.99483, -14.99903, -14.99967, -14.99903, 
    -14.99483, -14.98581, -14.97744, 0,
  0, -14.9994, -14.98064, -14.98906, -14.99483, -14.99644, -14.99483, 
    -14.98906, -14.98064, -14.9994, 0,
  0, -15, -14.99846, -14.98064, -14.98581, -14.98509, -14.98581, -14.98064, 
    -14.99846, -15, 0,
  0, 0, -15, -14.9994, -14.97744, -14.96799, -14.97744, -14.9994, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99865, -14.97534, -14.96512, -14.97534, -14.99865, -15, 0, 0,
  0, -15, -14.99625, -14.94263, -14.97022, -14.97184, -14.97022, -14.94263, 
    -14.99625, -15, 0,
  0, -14.99865, -14.94263, -14.97897, -14.98979, -14.99253, -14.98979, 
    -14.97897, -14.94263, -14.99865, 0,
  0, -14.97534, -14.97022, -14.98979, -14.99683, -14.99798, -14.99683, 
    -14.98979, -14.97022, -14.97534, 0,
  0, -14.96512, -14.97184, -14.99253, -14.99798, -14.99856, -14.99798, 
    -14.99253, -14.97184, -14.96512, 0,
  0, -14.97534, -14.97022, -14.98979, -14.99683, -14.99798, -14.99683, 
    -14.98979, -14.97022, -14.97534, 0,
  0, -14.99865, -14.94263, -14.97897, -14.98979, -14.99253, -14.98979, 
    -14.97897, -14.94263, -14.99865, 0,
  0, -15, -14.99625, -14.94263, -14.97022, -14.97184, -14.97022, -14.94263, 
    -14.99625, -15, 0,
  0, 0, -15, -14.99865, -14.97534, -14.96512, -14.97534, -14.99865, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99781, -14.97328, -14.96243, -14.97328, -14.99781, -15, 0, 0,
  0, -15, -14.99341, -14.84747, -14.9075, -14.9162, -14.9075, -14.84747, 
    -14.99341, -15, 0,
  0, -14.99781, -14.84747, -14.93055, -14.95609, -14.96239, -14.95609, 
    -14.93055, -14.84747, -14.99781, 0,
  0, -14.97328, -14.9075, -14.95609, -14.97254, -14.97591, -14.97254, 
    -14.95609, -14.9075, -14.97328, 0,
  0, -14.96243, -14.9162, -14.96239, -14.97591, -14.97832, -14.97591, 
    -14.96239, -14.9162, -14.96243, 0,
  0, -14.97328, -14.9075, -14.95609, -14.97254, -14.97591, -14.97254, 
    -14.95609, -14.9075, -14.97328, 0,
  0, -14.99781, -14.84747, -14.93055, -14.95609, -14.96239, -14.95609, 
    -14.93055, -14.84747, -14.99781, 0,
  0, -15, -14.99341, -14.84747, -14.9075, -14.9162, -14.9075, -14.84747, 
    -14.99341, -15, 0,
  0, 0, -15, -14.99781, -14.97328, -14.96243, -14.97328, -14.99781, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99837, -14.97183, -14.96027, -14.97183, -14.99837, -15, 0, 0,
  0, -15, -14.99452, -14.67498, -14.71689, -14.72601, -14.71689, -14.67498, 
    -14.99452, -15, 0,
  0, -14.99837, -14.67498, -14.74268, -14.77814, -14.78795, -14.77814, 
    -14.74268, -14.67498, -14.99837, 0,
  0, -14.97183, -14.71689, -14.77814, -14.80483, -14.81124, -14.80483, 
    -14.77814, -14.71689, -14.97183, 0,
  0, -14.96027, -14.72601, -14.78795, -14.81124, -14.8165, -14.81124, 
    -14.78795, -14.72601, -14.96027, 0,
  0, -14.97183, -14.71689, -14.77814, -14.80483, -14.81124, -14.80483, 
    -14.77814, -14.71689, -14.97183, 0,
  0, -14.99837, -14.67498, -14.74268, -14.77814, -14.78795, -14.77814, 
    -14.74268, -14.67498, -14.99837, 0,
  0, -15, -14.99452, -14.67498, -14.71689, -14.72601, -14.71689, -14.67498, 
    -14.99452, -15, 0,
  0, 0, -15, -14.99837, -14.97183, -14.96027, -14.97183, -14.99837, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -14.97207, -14.96025, -14.97207, -15, -15, -15, -15,
  -15, -15, -15, -14.54677, -14.51873, -14.50966, -14.51873, -14.54677, -15, 
    -15, -15,
  -15, -15, -14.54677, -14.50978, -14.50106, -14.4976, -14.50106, -14.50978, 
    -14.54677, -15, -15,
  -15, -14.97207, -14.51873, -14.50106, -14.48895, -14.48321, -14.48895, 
    -14.50106, -14.51873, -14.97207, -15,
  -15, -14.96025, -14.50966, -14.4976, -14.48321, -14.47674, -14.48321, 
    -14.4976, -14.50966, -14.96025, -15,
  -15, -14.97207, -14.51873, -14.50106, -14.48895, -14.48321, -14.48895, 
    -14.50106, -14.51873, -14.97207, -15,
  -15, -15, -14.54677, -14.50978, -14.50106, -14.4976, -14.50106, -14.50978, 
    -14.54677, -15, -15,
  -15, -15, -15, -14.54677, -14.51873, -14.50966, -14.51873, -14.54677, -15, 
    -15, -15,
  -15, -15, -15, -15, -14.97207, -14.96025, -14.97207, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99999, -14.99647, -14.99498, -14.99647, -14.99999, -15, 0, 0,
  0, -15, -14.99997, -14.99975, -14.99971, -14.99955, -14.99971, -14.99975, 
    -14.99997, -15, 0,
  0, -14.99999, -14.99975, -14.99978, -14.9997, -14.99968, -14.9997, 
    -14.99978, -14.99975, -14.99999, 0,
  0, -14.99647, -14.99971, -14.9997, -14.99985, -14.99994, -14.99985, 
    -14.9997, -14.99971, -14.99647, 0,
  0, -14.99498, -14.99955, -14.99968, -14.99994, -14.99999, -14.99994, 
    -14.99968, -14.99955, -14.99498, 0,
  0, -14.99647, -14.99971, -14.9997, -14.99985, -14.99994, -14.99985, 
    -14.9997, -14.99971, -14.99647, 0,
  0, -14.99999, -14.99975, -14.99978, -14.9997, -14.99968, -14.9997, 
    -14.99978, -14.99975, -14.99999, 0,
  0, -15, -14.99997, -14.99975, -14.99971, -14.99955, -14.99971, -14.99975, 
    -14.99997, -15, 0,
  0, 0, -15, -14.99999, -14.99647, -14.99498, -14.99647, -14.99999, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99997, -14.9904, -14.98636, -14.9904, -14.99997, -15, 0, 0,
  0, -15, -14.99993, -14.99934, -14.99926, -14.99903, -14.99926, -14.99934, 
    -14.99993, -15, 0,
  0, -14.99997, -14.99934, -14.99941, -14.9995, -14.99954, -14.9995, 
    -14.99941, -14.99934, -14.99997, 0,
  0, -14.9904, -14.99926, -14.9995, -14.9998, -14.99992, -14.9998, -14.9995, 
    -14.99926, -14.9904, 0,
  0, -14.98636, -14.99903, -14.99954, -14.99992, -15, -14.99992, -14.99954, 
    -14.99903, -14.98636, 0,
  0, -14.9904, -14.99926, -14.9995, -14.9998, -14.99992, -14.9998, -14.9995, 
    -14.99926, -14.9904, 0,
  0, -14.99997, -14.99934, -14.99941, -14.9995, -14.99954, -14.9995, 
    -14.99941, -14.99934, -14.99997, 0,
  0, -15, -14.99993, -14.99934, -14.99926, -14.99903, -14.99926, -14.99934, 
    -14.99993, -15, 0,
  0, 0, -15, -14.99997, -14.9904, -14.98636, -14.9904, -14.99997, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99991, -14.98569, -14.97974, -14.98569, -14.99991, -15, 0, 0,
  0, -15, -14.99981, -14.99811, -14.99772, -14.99741, -14.99772, -14.99811, 
    -14.99981, -15, 0,
  0, -14.99991, -14.99811, -14.99812, -14.99892, -14.99915, -14.99892, 
    -14.99812, -14.99811, -14.99991, 0,
  0, -14.98569, -14.99772, -14.99892, -14.9997, -14.99989, -14.9997, 
    -14.99892, -14.99772, -14.98569, 0,
  0, -14.97974, -14.99741, -14.99915, -14.99989, -15, -14.99989, -14.99915, 
    -14.99741, -14.97974, 0,
  0, -14.98569, -14.99772, -14.99892, -14.9997, -14.99989, -14.9997, 
    -14.99892, -14.99772, -14.98569, 0,
  0, -14.99991, -14.99811, -14.99812, -14.99892, -14.99915, -14.99892, 
    -14.99812, -14.99811, -14.99991, 0,
  0, -15, -14.99981, -14.99811, -14.99772, -14.99741, -14.99772, -14.99811, 
    -14.99981, -15, 0,
  0, 0, -15, -14.99991, -14.98569, -14.97974, -14.98569, -14.99991, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99983, -14.98194, -14.97443, -14.98194, -14.99983, -15, 0, 0,
  0, -15, -14.99963, -14.99574, -14.99479, -14.99429, -14.99479, -14.99574, 
    -14.99963, -15, 0,
  0, -14.99983, -14.99574, -14.99564, -14.9978, -14.99842, -14.9978, 
    -14.99564, -14.99574, -14.99983, 0,
  0, -14.98194, -14.99479, -14.9978, -14.99953, -14.99985, -14.99953, 
    -14.9978, -14.99479, -14.98194, 0,
  0, -14.97443, -14.99429, -14.99842, -14.99985, -15, -14.99985, -14.99842, 
    -14.99429, -14.97443, 0,
  0, -14.98194, -14.99479, -14.9978, -14.99953, -14.99985, -14.99953, 
    -14.9978, -14.99479, -14.98194, 0,
  0, -14.99983, -14.99574, -14.99564, -14.9978, -14.99842, -14.9978, 
    -14.99564, -14.99574, -14.99983, 0,
  0, -15, -14.99963, -14.99574, -14.99479, -14.99429, -14.99479, -14.99574, 
    -14.99963, -15, 0,
  0, 0, -15, -14.99983, -14.98194, -14.97443, -14.98194, -14.99983, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99969, -14.97893, -14.97014, -14.97893, -14.99969, -15, 0, 0,
  0, -15, -14.99928, -14.99083, -14.99062, -14.98987, -14.99062, -14.99083, 
    -14.99928, -15, 0,
  0, -14.99969, -14.99083, -14.99216, -14.99621, -14.99737, -14.99621, 
    -14.99216, -14.99083, -14.99969, 0,
  0, -14.97893, -14.99062, -14.99621, -14.99928, -14.99978, -14.99928, 
    -14.99621, -14.99062, -14.97893, 0,
  0, -14.97014, -14.98987, -14.99737, -14.99978, -15, -14.99978, -14.99737, 
    -14.98987, -14.97014, 0,
  0, -14.97893, -14.99062, -14.99621, -14.99928, -14.99978, -14.99928, 
    -14.99621, -14.99062, -14.97893, 0,
  0, -14.99969, -14.99083, -14.99216, -14.99621, -14.99737, -14.99621, 
    -14.99216, -14.99083, -14.99969, 0,
  0, -15, -14.99928, -14.99083, -14.99062, -14.98987, -14.99062, -14.99083, 
    -14.99928, -15, 0,
  0, 0, -15, -14.99969, -14.97893, -14.97014, -14.97893, -14.99969, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99923, -14.97643, -14.96664, -14.97643, -14.99923, -15, 0, 0,
  0, -15, -14.99812, -14.97587, -14.98409, -14.98359, -14.98409, -14.97587, 
    -14.99812, -15, 0,
  0, -14.99923, -14.97587, -14.98734, -14.99405, -14.9959, -14.99405, 
    -14.98734, -14.97587, -14.99923, 0,
  0, -14.97643, -14.98409, -14.99405, -14.99885, -14.9996, -14.99885, 
    -14.99405, -14.98409, -14.97643, 0,
  0, -14.96664, -14.98359, -14.9959, -14.9996, -14.99991, -14.9996, -14.9959, 
    -14.98359, -14.96664, 0,
  0, -14.97643, -14.98409, -14.99405, -14.99885, -14.9996, -14.99885, 
    -14.99405, -14.98409, -14.97643, 0,
  0, -14.99923, -14.97587, -14.98734, -14.99405, -14.9959, -14.99405, 
    -14.98734, -14.97587, -14.99923, 0,
  0, -15, -14.99812, -14.97587, -14.98409, -14.98359, -14.98409, -14.97587, 
    -14.99812, -15, 0,
  0, 0, -15, -14.99923, -14.97643, -14.96664, -14.97643, -14.99923, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.9984, -14.97421, -14.96369, -14.97421, -14.9984, -15, 0, 0,
  0, -15, -14.99588, -14.93004, -14.96479, -14.96736, -14.96479, -14.93004, 
    -14.99588, -15, 0,
  0, -14.9984, -14.93004, -14.97464, -14.98759, -14.99084, -14.98759, 
    -14.97464, -14.93004, -14.9984, 0,
  0, -14.97421, -14.96479, -14.98759, -14.99591, -14.99729, -14.99591, 
    -14.98759, -14.96479, -14.97421, 0,
  0, -14.96369, -14.96736, -14.99084, -14.99729, -14.998, -14.99729, 
    -14.99084, -14.96736, -14.96369, 0,
  0, -14.97421, -14.96479, -14.98759, -14.99591, -14.99729, -14.99591, 
    -14.98759, -14.96479, -14.97421, 0,
  0, -14.9984, -14.93004, -14.97464, -14.98759, -14.99084, -14.98759, 
    -14.97464, -14.93004, -14.9984, 0,
  0, -15, -14.99588, -14.93004, -14.96479, -14.96736, -14.96479, -14.93004, 
    -14.99588, -15, 0,
  0, 0, -15, -14.9984, -14.97421, -14.96369, -14.97421, -14.9984, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99756, -14.97203, -14.96081, -14.97203, -14.99756, -15, 0, 0,
  0, -15, -14.99329, -14.82399, -14.89138, -14.90177, -14.89138, -14.82399, 
    -14.99329, -15, 0,
  0, -14.99756, -14.82399, -14.91676, -14.9466, -14.95401, -14.9466, 
    -14.91676, -14.82399, -14.99756, 0,
  0, -14.97203, -14.89138, -14.9466, -14.96597, -14.97, -14.96597, -14.9466, 
    -14.89138, -14.97203, 0,
  0, -14.96081, -14.90177, -14.95401, -14.97, -14.97293, -14.97, -14.95401, 
    -14.90177, -14.96081, 0,
  0, -14.97203, -14.89138, -14.9466, -14.96597, -14.97, -14.96597, -14.9466, 
    -14.89138, -14.97203, 0,
  0, -14.99756, -14.82399, -14.91676, -14.9466, -14.95401, -14.9466, 
    -14.91676, -14.82399, -14.99756, 0,
  0, -15, -14.99329, -14.82399, -14.89138, -14.90177, -14.89138, -14.82399, 
    -14.99329, -15, 0,
  0, 0, -15, -14.99756, -14.97203, -14.96081, -14.97203, -14.99756, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99829, -14.97057, -14.9586, -14.97057, -14.99829, -15, 0, 0,
  0, -15, -14.99481, -14.64408, -14.68719, -14.69682, -14.68719, -14.64408, 
    -14.99481, -15, 0,
  0, -14.99829, -14.64408, -14.71307, -14.75152, -14.76225, -14.75152, 
    -14.71307, -14.64408, -14.99829, 0,
  0, -14.97057, -14.68719, -14.75152, -14.78076, -14.78779, -14.78076, 
    -14.75152, -14.68719, -14.97057, 0,
  0, -14.9586, -14.69682, -14.76225, -14.78779, -14.79355, -14.78779, 
    -14.76225, -14.69682, -14.9586, 0,
  0, -14.97057, -14.68719, -14.75152, -14.78076, -14.78779, -14.78076, 
    -14.75152, -14.68719, -14.97057, 0,
  0, -14.99829, -14.64408, -14.71307, -14.75152, -14.76225, -14.75152, 
    -14.71307, -14.64408, -14.99829, 0,
  0, -15, -14.99481, -14.64408, -14.68719, -14.69682, -14.68719, -14.64408, 
    -14.99481, -15, 0,
  0, 0, -15, -14.99829, -14.97057, -14.9586, -14.97057, -14.99829, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -14.97086, -14.95862, -14.97086, -15, -15, -15, -15,
  -15, -15, -15, -14.51575, -14.48891, -14.48036, -14.48891, -14.51575, -15, 
    -15, -15,
  -15, -15, -14.51575, -14.48022, -14.47459, -14.47206, -14.47459, -14.48022, 
    -14.51575, -15, -15,
  -15, -14.97086, -14.48891, -14.47459, -14.46499, -14.45983, -14.46499, 
    -14.47459, -14.48891, -14.97086, -15,
  -15, -14.95862, -14.48036, -14.47206, -14.45983, -14.45381, -14.45983, 
    -14.47206, -14.48036, -14.95862, -15,
  -15, -14.97086, -14.48891, -14.47459, -14.46499, -14.45983, -14.46499, 
    -14.47459, -14.48891, -14.97086, -15,
  -15, -15, -14.51575, -14.48022, -14.47459, -14.47206, -14.47459, -14.48022, 
    -14.51575, -15, -15,
  -15, -15, -15, -14.51575, -14.48891, -14.48036, -14.48891, -14.51575, -15, 
    -15, -15,
  -15, -15, -15, -15, -14.97086, -14.95862, -14.97086, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99998, -14.99631, -14.99478, -14.99631, -14.99998, -15, 0, 0,
  0, -15, -14.99997, -14.99972, -14.99969, -14.99953, -14.99969, -14.99972, 
    -14.99997, -15, 0,
  0, -14.99998, -14.99972, -14.99976, -14.99966, -14.99965, -14.99966, 
    -14.99976, -14.99972, -14.99998, 0,
  0, -14.99631, -14.99969, -14.99966, -14.99983, -14.99993, -14.99983, 
    -14.99966, -14.99969, -14.99631, 0,
  0, -14.99478, -14.99953, -14.99965, -14.99993, -14.99999, -14.99993, 
    -14.99965, -14.99953, -14.99478, 0,
  0, -14.99631, -14.99969, -14.99966, -14.99983, -14.99993, -14.99983, 
    -14.99966, -14.99969, -14.99631, 0,
  0, -14.99998, -14.99972, -14.99976, -14.99966, -14.99965, -14.99966, 
    -14.99976, -14.99972, -14.99998, 0,
  0, -15, -14.99997, -14.99972, -14.99969, -14.99953, -14.99969, -14.99972, 
    -14.99997, -15, 0,
  0, 0, -15, -14.99998, -14.99631, -14.99478, -14.99631, -14.99998, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99996, -14.98998, -14.9858, -14.98998, -14.99996, -15, 0, 0,
  0, -15, -14.99993, -14.99926, -14.99919, -14.99897, -14.99919, -14.99926, 
    -14.99993, -15, 0,
  0, -14.99996, -14.99926, -14.99933, -14.99944, -14.99949, -14.99944, 
    -14.99933, -14.99926, -14.99996, 0,
  0, -14.98998, -14.99919, -14.99944, -14.99978, -14.99991, -14.99978, 
    -14.99944, -14.99919, -14.98998, 0,
  0, -14.9858, -14.99897, -14.99949, -14.99991, -15, -14.99991, -14.99949, 
    -14.99897, -14.9858, 0,
  0, -14.98998, -14.99919, -14.99944, -14.99978, -14.99991, -14.99978, 
    -14.99944, -14.99919, -14.98998, 0,
  0, -14.99996, -14.99926, -14.99933, -14.99944, -14.99949, -14.99944, 
    -14.99933, -14.99926, -14.99996, 0,
  0, -15, -14.99993, -14.99926, -14.99919, -14.99897, -14.99919, -14.99926, 
    -14.99993, -15, 0,
  0, 0, -15, -14.99996, -14.98998, -14.9858, -14.98998, -14.99996, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99991, -14.98507, -14.97891, -14.98507, -14.99991, -15, 0, 0,
  0, -15, -14.99981, -14.99788, -14.99753, -14.99722, -14.99753, -14.99788, 
    -14.99981, -15, 0,
  0, -14.99991, -14.99788, -14.99789, -14.99879, -14.99905, -14.99879, 
    -14.99789, -14.99788, -14.99991, 0,
  0, -14.98507, -14.99753, -14.99879, -14.99966, -14.99988, -14.99966, 
    -14.99879, -14.99753, -14.98507, 0,
  0, -14.97891, -14.99722, -14.99905, -14.99988, -15, -14.99988, -14.99905, 
    -14.99722, -14.97891, 0,
  0, -14.98507, -14.99753, -14.99879, -14.99966, -14.99988, -14.99966, 
    -14.99879, -14.99753, -14.98507, 0,
  0, -14.99991, -14.99788, -14.99789, -14.99879, -14.99905, -14.99879, 
    -14.99789, -14.99788, -14.99991, 0,
  0, -15, -14.99981, -14.99788, -14.99753, -14.99722, -14.99753, -14.99788, 
    -14.99981, -15, 0,
  0, 0, -15, -14.99991, -14.98507, -14.97891, -14.98507, -14.99991, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99982, -14.98116, -14.97339, -14.98116, -14.99982, -15, 0, 0,
  0, -15, -14.99961, -14.99516, -14.99436, -14.99387, -14.99436, -14.99516, 
    -14.99961, -15, 0,
  0, -14.99982, -14.99516, -14.9951, -14.99753, -14.99823, -14.99753, 
    -14.9951, -14.99516, -14.99982, 0,
  0, -14.98116, -14.99436, -14.99753, -14.99947, -14.99983, -14.99947, 
    -14.99753, -14.99436, -14.98116, 0,
  0, -14.97339, -14.99387, -14.99823, -14.99983, -15, -14.99983, -14.99823, 
    -14.99387, -14.97339, 0,
  0, -14.98116, -14.99436, -14.99753, -14.99947, -14.99983, -14.99947, 
    -14.99753, -14.99436, -14.98116, 0,
  0, -14.99982, -14.99516, -14.9951, -14.99753, -14.99823, -14.99753, 
    -14.9951, -14.99516, -14.99982, 0,
  0, -15, -14.99961, -14.99516, -14.99436, -14.99387, -14.99436, -14.99516, 
    -14.99961, -15, 0,
  0, 0, -15, -14.99982, -14.98116, -14.97339, -14.98116, -14.99982, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99964, -14.97802, -14.96892, -14.97802, -14.99964, -15, 0, 0,
  0, -15, -14.99921, -14.98914, -14.9898, -14.98909, -14.9898, -14.98914, 
    -14.99921, -15, 0,
  0, -14.99964, -14.98914, -14.99118, -14.99575, -14.99705, -14.99575, 
    -14.99118, -14.98914, -14.99964, 0,
  0, -14.97802, -14.9898, -14.99575, -14.99918, -14.99975, -14.99918, 
    -14.99575, -14.9898, -14.97802, 0,
  0, -14.96892, -14.98909, -14.99705, -14.99975, -15, -14.99975, -14.99705, 
    -14.98909, -14.96892, 0,
  0, -14.97802, -14.9898, -14.99575, -14.99918, -14.99975, -14.99918, 
    -14.99575, -14.9898, -14.97802, 0,
  0, -14.99964, -14.98914, -14.99118, -14.99575, -14.99705, -14.99575, 
    -14.99118, -14.98914, -14.99964, 0,
  0, -15, -14.99921, -14.98914, -14.9898, -14.98909, -14.9898, -14.98914, 
    -14.99921, -15, 0,
  0, 0, -15, -14.99964, -14.97802, -14.96892, -14.97802, -14.99964, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.9991, -14.97542, -14.96529, -14.97542, -14.9991, -15, 0, 0,
  0, -15, -14.99793, -14.97058, -14.98222, -14.98199, -14.98222, -14.97058, 
    -14.99793, -15, 0,
  0, -14.9991, -14.97058, -14.98555, -14.99323, -14.99533, -14.99323, 
    -14.98555, -14.97058, -14.9991, 0,
  0, -14.97542, -14.98222, -14.99323, -14.99866, -14.99951, -14.99866, 
    -14.99323, -14.98222, -14.97542, 0,
  0, -14.96529, -14.98199, -14.99533, -14.99951, -14.99988, -14.99951, 
    -14.99533, -14.98199, -14.96529, 0,
  0, -14.97542, -14.98222, -14.99323, -14.99866, -14.99951, -14.99866, 
    -14.99323, -14.98222, -14.97542, 0,
  0, -14.9991, -14.97058, -14.98555, -14.99323, -14.99533, -14.99323, 
    -14.98555, -14.97058, -14.9991, 0,
  0, -15, -14.99793, -14.97058, -14.98222, -14.98199, -14.98222, -14.97058, 
    -14.99793, -15, 0,
  0, 0, -15, -14.9991, -14.97542, -14.96529, -14.97542, -14.9991, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99817, -14.97307, -14.96219, -14.97307, -14.99817, -15, 0, 0,
  0, -15, -14.9956, -14.91692, -14.95888, -14.96247, -14.95888, -14.91692, 
    -14.9956, -15, 0,
  0, -14.99817, -14.91692, -14.96996, -14.98516, -14.98895, -14.98516, 
    -14.96996, -14.91692, -14.99817, 0,
  0, -14.97307, -14.95888, -14.98516, -14.99483, -14.99647, -14.99483, 
    -14.98516, -14.95888, -14.97307, 0,
  0, -14.96219, -14.96247, -14.98895, -14.99647, -14.99734, -14.99647, 
    -14.98895, -14.96247, -14.96219, 0,
  0, -14.97307, -14.95888, -14.98516, -14.99483, -14.99647, -14.99483, 
    -14.98516, -14.95888, -14.97307, 0,
  0, -14.99817, -14.91692, -14.96996, -14.98516, -14.98895, -14.98516, 
    -14.96996, -14.91692, -14.99817, 0,
  0, -15, -14.9956, -14.91692, -14.95888, -14.96247, -14.95888, -14.91692, 
    -14.9956, -15, 0,
  0, 0, -15, -14.99817, -14.97307, -14.96219, -14.97307, -14.99817, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99734, -14.97078, -14.95918, -14.97078, -14.99734, -15, 0, 0,
  0, -15, -14.99321, -14.80103, -14.87498, -14.88696, -14.87498, -14.80103, 
    -14.99321, -15, 0,
  0, -14.99734, -14.80103, -14.90252, -14.93661, -14.94514, -14.93661, 
    -14.90252, -14.80103, -14.99734, 0,
  0, -14.97078, -14.87498, -14.93661, -14.95895, -14.96366, -14.95895, 
    -14.93661, -14.87498, -14.97078, 0,
  0, -14.95918, -14.88696, -14.94514, -14.96366, -14.96712, -14.96366, 
    -14.94514, -14.88696, -14.95918, 0,
  0, -14.97078, -14.87498, -14.93661, -14.95895, -14.96366, -14.95895, 
    -14.93661, -14.87498, -14.97078, 0,
  0, -14.99734, -14.80103, -14.90252, -14.93661, -14.94514, -14.93661, 
    -14.90252, -14.80103, -14.99734, 0,
  0, -15, -14.99321, -14.80103, -14.87498, -14.88696, -14.87498, -14.80103, 
    -14.99321, -15, 0,
  0, 0, -15, -14.99734, -14.97078, -14.95918, -14.97078, -14.99734, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -15, -14.99821, -14.96931, -14.95693, -14.96931, -14.99821, -15, 0, 0,
  0, -15, -14.99505, -14.61492, -14.65891, -14.66894, -14.65891, -14.61492, 
    -14.99505, -15, 0,
  0, -14.99821, -14.61492, -14.68469, -14.72585, -14.73743, -14.72585, 
    -14.68469, -14.61492, -14.99821, 0,
  0, -14.96931, -14.65891, -14.72585, -14.75744, -14.76506, -14.75744, 
    -14.72585, -14.65891, -14.96931, 0,
  0, -14.95693, -14.66894, -14.73743, -14.76506, -14.77127, -14.76506, 
    -14.73743, -14.66894, -14.95693, 0,
  0, -14.96931, -14.65891, -14.72585, -14.75744, -14.76506, -14.75744, 
    -14.72585, -14.65891, -14.96931, 0,
  0, -14.99821, -14.61492, -14.68469, -14.72585, -14.73743, -14.72585, 
    -14.68469, -14.61492, -14.99821, 0,
  0, -15, -14.99505, -14.61492, -14.65891, -14.66894, -14.65891, -14.61492, 
    -14.99505, -15, 0,
  0, 0, -15, -14.99821, -14.96931, -14.95693, -14.96931, -14.99821, -15, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -14.96965, -14.95699, -14.96965, -15, -15, -15, -15,
  -15, -15, -15, -14.48647, -14.46052, -14.45237, -14.46052, -14.48647, -15, 
    -15, -15,
  -15, -15, -14.48647, -14.45189, -14.44908, -14.4474, -14.44908, -14.45189, 
    -14.48647, -15, -15,
  -15, -14.96965, -14.46052, -14.44908, -14.44179, -14.43715, -14.44179, 
    -14.44908, -14.46052, -14.96965, -15,
  -15, -14.95699, -14.45237, -14.4474, -14.43715, -14.43154, -14.43715, 
    -14.4474, -14.45237, -14.95699, -15,
  -15, -14.96965, -14.46052, -14.44908, -14.44179, -14.43715, -14.44179, 
    -14.44908, -14.46052, -14.96965, -15,
  -15, -15, -14.48647, -14.45189, -14.44908, -14.4474, -14.44908, -14.45189, 
    -14.48647, -15, -15,
  -15, -15, -15, -14.48647, -14.46052, -14.45237, -14.46052, -14.48647, -15, 
    -15, -15,
  -15, -15, -15, -15, -14.96965, -14.95699, -14.96965, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -15, -14.99999, -14.99615, -14.99458, -14.99615, -14.99999, -15, 
    -15, 0,
  0, -15, -14.99702, -14.99969, -14.99967, -14.99952, -14.99967, -14.99969, 
    -14.99702, -15, 0,
  0, -14.99999, -14.99969, -14.99974, -14.99963, -14.99961, -14.99963, 
    -14.99974, -14.99969, -14.99999, 0,
  0, -14.99615, -14.99967, -14.99963, -14.99982, -14.99992, -14.99982, 
    -14.99963, -14.99967, -14.99615, 0,
  0, -14.99458, -14.99952, -14.99961, -14.99992, -14.99999, -14.99992, 
    -14.99961, -14.99952, -14.99458, 0,
  0, -14.99615, -14.99967, -14.99963, -14.99982, -14.99992, -14.99982, 
    -14.99963, -14.99967, -14.99615, 0,
  0, -14.99999, -14.99969, -14.99974, -14.99963, -14.99961, -14.99963, 
    -14.99974, -14.99969, -14.99999, 0,
  0, -15, -14.99702, -14.99969, -14.99967, -14.99952, -14.99967, -14.99969, 
    -14.99702, -15, 0,
  0, -15, -15, -14.99999, -14.99615, -14.99458, -14.99615, -14.99999, -15, 
    -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -14.99999, -14.99999, -14.98953, -14.98526, -14.98953, -14.99999, 
    -14.99999, -15, 0,
  0, -14.99999, -14.99188, -14.9992, -14.99913, -14.99891, -14.99913, 
    -14.9992, -14.99188, -14.99999, 0,
  0, -14.99999, -14.9992, -14.99928, -14.99939, -14.99944, -14.99939, 
    -14.99928, -14.9992, -14.99999, 0,
  0, -14.98953, -14.99913, -14.99939, -14.99976, -14.9999, -14.99976, 
    -14.99939, -14.99913, -14.98953, 0,
  0, -14.98526, -14.99891, -14.99944, -14.9999, -14.99999, -14.9999, 
    -14.99944, -14.99891, -14.98526, 0,
  0, -14.98953, -14.99913, -14.99939, -14.99976, -14.9999, -14.99976, 
    -14.99939, -14.99913, -14.98953, 0,
  0, -14.99999, -14.9992, -14.99928, -14.99939, -14.99944, -14.99939, 
    -14.99928, -14.9992, -14.99999, 0,
  0, -14.99999, -14.99188, -14.9992, -14.99913, -14.99891, -14.99913, 
    -14.9992, -14.99188, -14.99999, 0,
  0, -15, -14.99999, -14.99999, -14.98953, -14.98526, -14.98953, -14.99999, 
    -14.99999, -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -14.99999, -14.99997, -14.98441, -14.97809, -14.98441, -14.99997, 
    -14.99999, -15, 0,
  0, -14.99999, -14.98794, -14.99773, -14.99734, -14.99703, -14.99734, 
    -14.99773, -14.98794, -14.99999, 0,
  0, -14.99997, -14.99773, -14.99771, -14.99866, -14.99896, -14.99866, 
    -14.99771, -14.99773, -14.99997, 0,
  0, -14.98441, -14.99734, -14.99866, -14.99963, -14.99986, -14.99963, 
    -14.99866, -14.99734, -14.98441, 0,
  0, -14.97809, -14.99703, -14.99896, -14.99986, -15, -14.99986, -14.99896, 
    -14.99703, -14.97809, 0,
  0, -14.98441, -14.99734, -14.99866, -14.99963, -14.99986, -14.99963, 
    -14.99866, -14.99734, -14.98441, 0,
  0, -14.99997, -14.99773, -14.99771, -14.99866, -14.99896, -14.99866, 
    -14.99771, -14.99773, -14.99997, 0,
  0, -14.99999, -14.98794, -14.99773, -14.99734, -14.99703, -14.99734, 
    -14.99773, -14.98794, -14.99999, 0,
  0, -15, -14.99999, -14.99997, -14.98441, -14.97809, -14.98441, -14.99997, 
    -14.99999, -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -14.99999, -14.99993, -14.98035, -14.97235, -14.98035, -14.99993, 
    -14.99999, -15, 0,
  0, -14.99999, -14.98484, -14.99473, -14.99394, -14.99344, -14.99394, 
    -14.99473, -14.98484, -14.99999, 0,
  0, -14.99993, -14.99473, -14.9947, -14.99727, -14.99805, -14.99727, 
    -14.9947, -14.99473, -14.99993, 0,
  0, -14.98035, -14.99394, -14.99727, -14.99941, -14.99981, -14.99941, 
    -14.99727, -14.99394, -14.98035, 0,
  0, -14.97235, -14.99344, -14.99805, -14.99981, -15, -14.99981, -14.99805, 
    -14.99344, -14.97235, 0,
  0, -14.98035, -14.99394, -14.99727, -14.99941, -14.99981, -14.99941, 
    -14.99727, -14.99394, -14.98035, 0,
  0, -14.99993, -14.99473, -14.9947, -14.99727, -14.99805, -14.99727, 
    -14.9947, -14.99473, -14.99993, 0,
  0, -14.99999, -14.98484, -14.99473, -14.99394, -14.99344, -14.99394, 
    -14.99473, -14.98484, -14.99999, 0,
  0, -15, -14.99999, -14.99993, -14.98035, -14.97235, -14.98035, -14.99993, 
    -14.99999, -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -14.99999, -14.9998, -14.97709, -14.96772, -14.97709, -14.9998, 
    -14.99999, -15, 0,
  0, -14.99999, -14.9823, -14.98759, -14.98898, -14.98829, -14.98898, 
    -14.98759, -14.9823, -14.99999, 0,
  0, -14.9998, -14.98759, -14.99043, -14.99529, -14.99673, -14.99529, 
    -14.99043, -14.98759, -14.9998, 0,
  0, -14.97709, -14.98898, -14.99529, -14.99909, -14.99972, -14.99909, 
    -14.99529, -14.98898, -14.97709, 0,
  0, -14.96772, -14.98829, -14.99673, -14.99972, -14.99999, -14.99972, 
    -14.99673, -14.98829, -14.96772, 0,
  0, -14.97709, -14.98898, -14.99529, -14.99909, -14.99972, -14.99909, 
    -14.99529, -14.98898, -14.97709, 0,
  0, -14.9998, -14.98759, -14.99043, -14.99529, -14.99673, -14.99529, 
    -14.99043, -14.98759, -14.9998, 0,
  0, -14.99999, -14.9823, -14.98759, -14.98898, -14.98829, -14.98898, 
    -14.98759, -14.9823, -14.99999, 0,
  0, -15, -14.99999, -14.9998, -14.97709, -14.96772, -14.97709, -14.9998, 
    -14.99999, -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -15, -14.99939, -14.97439, -14.96393, -14.97439, -14.99939, -15, 
    -15, 0,
  0, -15, -14.98005, -14.96531, -14.98025, -14.98027, -14.98025, -14.96531, 
    -14.98005, -15, 0,
  0, -14.99939, -14.96531, -14.98406, -14.99239, -14.99473, -14.99239, 
    -14.98406, -14.96531, -14.99939, 0,
  0, -14.97439, -14.98025, -14.99239, -14.99845, -14.99941, -14.99845, 
    -14.99239, -14.98025, -14.97439, 0,
  0, -14.96393, -14.98027, -14.99473, -14.99941, -14.99983, -14.99941, 
    -14.99473, -14.98027, -14.96393, 0,
  0, -14.97439, -14.98025, -14.99239, -14.99845, -14.99941, -14.99845, 
    -14.99239, -14.98025, -14.97439, 0,
  0, -14.99939, -14.96531, -14.98406, -14.99239, -14.99473, -14.99239, 
    -14.98406, -14.96531, -14.99939, 0,
  0, -15, -14.98005, -14.96531, -14.98025, -14.98027, -14.98025, -14.96531, 
    -14.98005, -15, 0,
  0, -15, -15, -14.99939, -14.97439, -14.96393, -14.97439, -14.99939, -15, 
    -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -15, -14.9988, -14.97194, -14.96066, -14.97194, -14.9988, -15, -15, 0,
  0, -15, -14.97781, -14.90411, -14.95259, -14.95718, -14.95259, -14.90411, 
    -14.97781, -15, 0,
  0, -14.9988, -14.90411, -14.96545, -14.98253, -14.98686, -14.98253, 
    -14.96545, -14.90411, -14.9988, 0,
  0, -14.97194, -14.95259, -14.98253, -14.99362, -14.99552, -14.99362, 
    -14.98253, -14.95259, -14.97194, 0,
  0, -14.96066, -14.95718, -14.98686, -14.99552, -14.99657, -14.99552, 
    -14.98686, -14.95718, -14.96066, 0,
  0, -14.97194, -14.95259, -14.98253, -14.99362, -14.99552, -14.99362, 
    -14.98253, -14.95259, -14.97194, 0,
  0, -14.9988, -14.90411, -14.96545, -14.98253, -14.98686, -14.98253, 
    -14.96545, -14.90411, -14.9988, 0,
  0, -15, -14.97781, -14.90411, -14.95259, -14.95718, -14.95259, -14.90411, 
    -14.97781, -15, 0,
  0, -15, -15, -14.9988, -14.97194, -14.96066, -14.97194, -14.9988, -15, -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -15, -14.99834, -14.96959, -14.95752, -14.96959, -14.99834, -15, 
    -15, 0,
  0, -15, -14.97594, -14.77949, -14.85847, -14.87185, -14.85847, -14.77949, 
    -14.97594, -15, 0,
  0, -14.99834, -14.77949, -14.88863, -14.92623, -14.93584, -14.92623, 
    -14.88863, -14.77949, -14.99834, 0,
  0, -14.96959, -14.85847, -14.92623, -14.95152, -14.95693, -14.95152, 
    -14.92623, -14.85847, -14.96959, 0,
  0, -14.95752, -14.87185, -14.93584, -14.95693, -14.96094, -14.95693, 
    -14.93584, -14.87185, -14.95752, 0,
  0, -14.96959, -14.85847, -14.92623, -14.95152, -14.95693, -14.95152, 
    -14.92623, -14.85847, -14.96959, 0,
  0, -14.99834, -14.77949, -14.88863, -14.92623, -14.93584, -14.92623, 
    -14.88863, -14.77949, -14.99834, 0,
  0, -15, -14.97594, -14.77949, -14.85847, -14.87185, -14.85847, -14.77949, 
    -14.97594, -15, 0,
  0, -15, -15, -14.99834, -14.96959, -14.95752, -14.96959, -14.99834, -15, 
    -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -15, -15, -14.99895, -14.96811, -14.95524, -14.96811, -14.99895, -15, 
    -15, 0,
  0, -15, -14.97532, -14.58826, -14.63196, -14.64219, -14.63196, -14.58826, 
    -14.97532, -15, 0,
  0, -14.99895, -14.58826, -14.6582, -14.70109, -14.71341, -14.70109, 
    -14.6582, -14.58826, -14.99895, 0,
  0, -14.96811, -14.63196, -14.70109, -14.73484, -14.74298, -14.73484, 
    -14.70109, -14.63196, -14.96811, 0,
  0, -14.95524, -14.64219, -14.71341, -14.74298, -14.74962, -14.74298, 
    -14.71341, -14.64219, -14.95524, 0,
  0, -14.96811, -14.63196, -14.70109, -14.73484, -14.74298, -14.73484, 
    -14.70109, -14.63196, -14.96811, 0,
  0, -14.99895, -14.58826, -14.6582, -14.70109, -14.71341, -14.70109, 
    -14.6582, -14.58826, -14.99895, 0,
  0, -15, -14.97532, -14.58826, -14.63196, -14.64219, -14.63196, -14.58826, 
    -14.97532, -15, 0,
  0, -15, -15, -14.99895, -14.96811, -14.95524, -14.96811, -14.99895, -15, 
    -15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -14.96843, -14.95534, -14.96843, -15, -15, -15, -15,
  -15, -15, -14.97576, -14.4597, -14.43346, -14.42552, -14.43346, -14.4597, 
    -14.97576, -15, -15,
  -15, -15, -14.4597, -14.42545, -14.42446, -14.42355, -14.42446, -14.42545, 
    -14.4597, -15, -15,
  -15, -14.96843, -14.43346, -14.42446, -14.4193, -14.41515, -14.4193, 
    -14.42446, -14.43346, -14.96843, -15,
  -15, -14.95534, -14.42552, -14.42355, -14.41515, -14.4099, -14.41515, 
    -14.42355, -14.42552, -14.95534, -15,
  -15, -14.96843, -14.43346, -14.42446, -14.4193, -14.41515, -14.4193, 
    -14.42446, -14.43346, -14.96843, -15,
  -15, -15, -14.4597, -14.42545, -14.42446, -14.42355, -14.42446, -14.42545, 
    -14.4597, -15, -15,
  -15, -15, -14.97576, -14.4597, -14.43346, -14.42552, -14.43346, -14.4597, 
    -14.97576, -15, -15,
  -15, -15, -15, -15, -14.96843, -14.95534, -14.96843, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 thk =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.1325216, 0.2058042, 0.2249885, 0.2058042, 0.1325216, 0, 0, 0,
  0, 0, 0.1325216, 0.2426609, 0.289271, 0.3032196, 0.289271, 0.2426609, 
    0.1325216, 0, 0,
  0, 0, 0.2058042, 0.289271, 0.3293495, 0.3416658, 0.3293495, 0.289271, 
    0.2058042, 0, 0,
  0, 0, 0.2249885, 0.3032196, 0.3416658, 0.3535534, 0.3416658, 0.3032196, 
    0.2249885, 0, 0,
  0, 0, 0.2058042, 0.289271, 0.3293495, 0.3416658, 0.3293495, 0.289271, 
    0.2058042, 0, 0,
  0, 0, 0.1325216, 0.2426609, 0.289271, 0.3032196, 0.289271, 0.2426609, 
    0.1325216, 0, 0,
  0, 0, 0, 0.1325216, 0.2058042, 0.2249885, 0.2058042, 0.1325216, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 3.201627e-05, 0.0002929367, 0.0005178058, 0.0002929367, 
    3.201627e-05, 0, 0, 0,
  0, 0, 5.686403e-05, 0.1326432, 0.2056712, 0.2245772, 0.2056712, 0.1326432, 
    5.686403e-05, 0, 0,
  0, 3.201627e-05, 0.1326432, 0.242601, 0.2890971, 0.3030184, 0.2890971, 
    0.242601, 0.1326432, 3.201627e-05, 0,
  0, 0.0002929367, 0.2056712, 0.2890971, 0.3292324, 0.3416044, 0.3292324, 
    0.2890971, 0.2056712, 0.0002929367, 0,
  0, 0.0005178058, 0.2245772, 0.3030184, 0.3416044, 0.3535409, 0.3416044, 
    0.3030184, 0.2245772, 0.0005178058, 0,
  0, 0.0002929367, 0.2056712, 0.2890971, 0.3292324, 0.3416044, 0.3292324, 
    0.2890971, 0.2056712, 0.0002929367, 0,
  0, 3.201627e-05, 0.1326432, 0.242601, 0.2890971, 0.3030184, 0.2890971, 
    0.242601, 0.1326432, 3.201627e-05, 0,
  0, 0, 5.686403e-05, 0.1326432, 0.2056712, 0.2245772, 0.2056712, 0.1326432, 
    5.686403e-05, 0, 0,
  0, 0, 0, 3.201627e-05, 0.0002929367, 0.0005178058, 0.0002929367, 
    3.201627e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3.499507e-10, 6.994776e-05, 0.0004022547, 0.0006260089, 0.0004022547, 
    6.994776e-05, 3.499507e-10, 0, 0,
  0, 3.499507e-10, 0.0001142617, 0.1327566, 0.205702, 0.2246232, 0.205702, 
    0.1327566, 0.0001142617, 3.499507e-10, 0,
  0, 6.994776e-05, 0.1327566, 0.2425436, 0.2889217, 0.302815, 0.2889217, 
    0.2425436, 0.1327566, 6.994776e-05, 0,
  0, 0.0004022547, 0.205702, 0.2889217, 0.3291154, 0.3415415, 0.3291154, 
    0.2889217, 0.205702, 0.0004022547, 0,
  0, 0.0006260089, 0.2246232, 0.302815, 0.3415415, 0.3535296, 0.3415415, 
    0.302815, 0.2246232, 0.0006260089, 0,
  0, 0.0004022547, 0.205702, 0.2889217, 0.3291154, 0.3415415, 0.3291154, 
    0.2889217, 0.205702, 0.0004022547, 0,
  0, 6.994776e-05, 0.1327566, 0.2425436, 0.2889217, 0.302815, 0.2889217, 
    0.2425436, 0.1327566, 6.994776e-05, 0,
  0, 3.499507e-10, 0.0001142617, 0.1327566, 0.205702, 0.2246232, 0.205702, 
    0.1327566, 0.0001142617, 3.499507e-10, 0,
  0, 0, 3.499507e-10, 6.994776e-05, 0.0004022547, 0.0006260089, 0.0004022547, 
    6.994776e-05, 3.499507e-10, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.146815e-09, 0.0001080381, 0.0005117886, 0.0007343993, 0.0005117886, 
    0.0001080381, 1.146815e-09, 0, 0,
  0, 1.146815e-09, 0.0001718189, 0.1328695, 0.2057316, 0.224668, 0.2057316, 
    0.1328695, 0.0001718189, 1.146815e-09, 0,
  0, 0.0001080381, 0.1328695, 0.2424858, 0.2887474, 0.3026132, 0.2887474, 
    0.2424858, 0.1328695, 0.0001080381, 0,
  0, 0.0005117886, 0.2057316, 0.2887474, 0.3289987, 0.3414782, 0.3289987, 
    0.2887474, 0.2057316, 0.0005117886, 0,
  0, 0.0007343993, 0.224668, 0.3026132, 0.3414782, 0.3535181, 0.3414782, 
    0.3026132, 0.224668, 0.0007343993, 0,
  0, 0.0005117886, 0.2057316, 0.2887474, 0.3289987, 0.3414782, 0.3289987, 
    0.2887474, 0.2057316, 0.0005117886, 0,
  0, 0.0001080381, 0.1328695, 0.2424858, 0.2887474, 0.3026132, 0.2887474, 
    0.2424858, 0.1328695, 0.0001080381, 0,
  0, 1.146815e-09, 0.0001718189, 0.1328695, 0.2057316, 0.224668, 0.2057316, 
    0.1328695, 0.0001718189, 1.146815e-09, 0,
  0, 0, 1.146815e-09, 0.0001080381, 0.0005117886, 0.0007343993, 0.0005117886, 
    0.0001080381, 1.146815e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3.71059e-09, 0.0001152924, 0.0005366366, 0.0007680521, 0.0005366366, 
    0.0001152924, 3.71059e-09, 0, 0,
  0, 3.71059e-09, 0.0002283403, 0.1329929, 0.2058461, 0.2247803, 0.2058461, 
    0.1329929, 0.0002283403, 3.71059e-09, 0,
  0, 0.0001152924, 0.1329929, 0.2424286, 0.2885876, 0.3024359, 0.2885876, 
    0.2424286, 0.1329929, 0.0001152924, 0,
  0, 0.0005366366, 0.2058461, 0.2885876, 0.3288787, 0.3414127, 0.3288787, 
    0.2885876, 0.2058461, 0.0005366366, 0,
  0, 0.0007680521, 0.2247803, 0.3024359, 0.3414127, 0.353507, 0.3414127, 
    0.3024359, 0.2247803, 0.0007680521, 0,
  0, 0.0005366366, 0.2058461, 0.2885876, 0.3288787, 0.3414127, 0.3288787, 
    0.2885876, 0.2058461, 0.0005366366, 0,
  0, 0.0001152924, 0.1329929, 0.2424286, 0.2885876, 0.3024359, 0.2885876, 
    0.2424286, 0.1329929, 0.0001152924, 0,
  0, 3.71059e-09, 0.0002283403, 0.1329929, 0.2058461, 0.2247803, 0.2058461, 
    0.1329929, 0.0002283403, 3.71059e-09, 0,
  0, 0, 3.71059e-09, 0.0001152924, 0.0005366366, 0.0007680521, 0.0005366366, 
    0.0001152924, 3.71059e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 7.089051e-09, 0.000122646, 0.0005616767, 0.0008019177, 0.0005616767, 
    0.000122646, 7.089051e-09, 0, 0,
  0, 7.089051e-09, 0.0002850269, 0.1331159, 0.2059595, 0.2248914, 0.2059595, 
    0.1331159, 0.0002850269, 7.089051e-09, 0,
  0, 0.000122646, 0.1331159, 0.2423711, 0.2884287, 0.30226, 0.2884287, 
    0.2423711, 0.1331159, 0.000122646, 0,
  0, 0.0005616767, 0.2059595, 0.2884287, 0.328759, 0.3413469, 0.328759, 
    0.2884287, 0.2059595, 0.0005616767, 0,
  0, 0.0008019177, 0.2248914, 0.30226, 0.3413469, 0.3534958, 0.3413469, 
    0.30226, 0.2248914, 0.0008019177, 0,
  0, 0.0005616767, 0.2059595, 0.2884287, 0.328759, 0.3413469, 0.328759, 
    0.2884287, 0.2059595, 0.0005616767, 0,
  0, 0.000122646, 0.1331159, 0.2423711, 0.2884287, 0.30226, 0.2884287, 
    0.2423711, 0.1331159, 0.000122646, 0,
  0, 7.089051e-09, 0.0002850269, 0.1331159, 0.2059595, 0.2248914, 0.2059595, 
    0.1331159, 0.0002850269, 7.089051e-09, 0,
  0, 0, 7.089051e-09, 0.000122646, 0.0005616767, 0.0008019177, 0.0005616767, 
    0.000122646, 7.089051e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.134039e-08, 0.0001300937, 0.0005868892, 0.0008359754, 0.0005868892, 
    0.0001300937, 1.134039e-08, 0, 0,
  0, 1.134039e-08, 0.0003418765, 0.1332385, 0.206072, 0.2250013, 0.206072, 
    0.1332385, 0.0003418765, 1.134039e-08, 0,
  0, 0.0001300937, 0.1332385, 0.2423133, 0.2882708, 0.3020855, 0.2882708, 
    0.2423133, 0.1332385, 0.0001300937, 0,
  0, 0.0005868892, 0.206072, 0.2882708, 0.3286397, 0.3412811, 0.3286397, 
    0.2882708, 0.206072, 0.0005868892, 0,
  0, 0.0008359754, 0.2250013, 0.3020855, 0.3412811, 0.3534843, 0.3412811, 
    0.3020855, 0.2250013, 0.0008359754, 0,
  0, 0.0005868892, 0.206072, 0.2882708, 0.3286397, 0.3412811, 0.3286397, 
    0.2882708, 0.206072, 0.0005868892, 0,
  0, 0.0001300937, 0.1332385, 0.2423133, 0.2882708, 0.3020855, 0.2882708, 
    0.2423133, 0.1332385, 0.0001300937, 0,
  0, 1.134039e-08, 0.0003418765, 0.1332385, 0.206072, 0.2250013, 0.206072, 
    0.1332385, 0.0003418765, 1.134039e-08, 0,
  0, 0, 1.134039e-08, 0.0001300937, 0.0005868892, 0.0008359754, 0.0005868892, 
    0.0001300937, 1.134039e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.651755e-08, 0.0001376354, 0.0006122729, 0.0008702234, 0.0006122729, 
    0.0001376354, 1.651755e-08, 0, 0,
  0, 1.651755e-08, 0.0003988868, 0.1333608, 0.2061835, 0.22511, 0.2061835, 
    0.1333608, 0.0003988868, 1.651755e-08, 0,
  0, 0.0001376354, 0.1333608, 0.2422552, 0.2881137, 0.3019123, 0.2881137, 
    0.2422552, 0.1333608, 0.0001376354, 0,
  0, 0.0006122729, 0.2061835, 0.2881137, 0.3285207, 0.341215, 0.3285207, 
    0.2881137, 0.2061835, 0.0006122729, 0,
  0, 0.0008702234, 0.22511, 0.3019123, 0.341215, 0.3534726, 0.341215, 
    0.3019123, 0.22511, 0.0008702234, 0,
  0, 0.0006122729, 0.2061835, 0.2881137, 0.3285207, 0.341215, 0.3285207, 
    0.2881137, 0.2061835, 0.0006122729, 0,
  0, 0.0001376354, 0.1333608, 0.2422552, 0.2881137, 0.3019123, 0.2881137, 
    0.2422552, 0.1333608, 0.0001376354, 0,
  0, 1.651755e-08, 0.0003988868, 0.1333608, 0.2061835, 0.22511, 0.2061835, 
    0.1333608, 0.0003988868, 1.651755e-08, 0,
  0, 0, 1.651755e-08, 0.0001376354, 0.0006122729, 0.0008702234, 0.0006122729, 
    0.0001376354, 1.651755e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 2.267689e-08, 0.0001452712, 0.0006378272, 0.0009046606, 0.0006378272, 
    0.0001452712, 2.267689e-08, 0, 0,
  0, 2.267689e-08, 0.0004560562, 0.1334826, 0.206294, 0.2252176, 0.206294, 
    0.1334826, 0.0004560562, 2.267689e-08, 0,
  0, 0.0001452712, 0.1334826, 0.2421968, 0.2879576, 0.3017404, 0.2879576, 
    0.2421968, 0.1334826, 0.0001452712, 0,
  0, 0.0006378272, 0.206294, 0.2879576, 0.3284021, 0.3411488, 0.3284021, 
    0.2879576, 0.206294, 0.0006378272, 0,
  0, 0.0009046606, 0.2252176, 0.3017404, 0.3411488, 0.3534607, 0.3411488, 
    0.3017404, 0.2252176, 0.0009046606, 0,
  0, 0.0006378272, 0.206294, 0.2879576, 0.3284021, 0.3411488, 0.3284021, 
    0.2879576, 0.206294, 0.0006378272, 0,
  0, 0.0001452712, 0.1334826, 0.2421968, 0.2879576, 0.3017404, 0.2879576, 
    0.2421968, 0.1334826, 0.0001452712, 0,
  0, 2.267689e-08, 0.0004560562, 0.1334826, 0.206294, 0.2252176, 0.206294, 
    0.1334826, 0.0004560562, 2.267689e-08, 0,
  0, 0, 2.267689e-08, 0.0001452712, 0.0006378272, 0.0009046606, 0.0006378272, 
    0.0001452712, 2.267689e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 2.987244e-08, 0.0001530009, 0.000663551, 0.0009392853, 0.000663551, 
    0.0001530009, 2.987244e-08, 0, 0,
  0, 2.987244e-08, 0.0005133827, 0.1336041, 0.2064035, 0.2253239, 0.2064035, 
    0.1336041, 0.0005133827, 2.987244e-08, 0,
  0, 0.0001530009, 0.1336041, 0.2421382, 0.2878024, 0.3015697, 0.2878024, 
    0.2421382, 0.1336041, 0.0001530009, 0,
  0, 0.000663551, 0.2064035, 0.2878024, 0.3282839, 0.3410824, 0.3282839, 
    0.2878024, 0.2064035, 0.000663551, 0,
  0, 0.0009392853, 0.2253239, 0.3015697, 0.3410824, 0.3534486, 0.3410824, 
    0.3015697, 0.2253239, 0.0009392853, 0,
  0, 0.000663551, 0.2064035, 0.2878024, 0.3282839, 0.3410824, 0.3282839, 
    0.2878024, 0.2064035, 0.000663551, 0,
  0, 0.0001530009, 0.1336041, 0.2421382, 0.2878024, 0.3015697, 0.2878024, 
    0.2421382, 0.1336041, 0.0001530009, 0,
  0, 2.987244e-08, 0.0005133827, 0.1336041, 0.2064035, 0.2253239, 0.2064035, 
    0.1336041, 0.0005133827, 2.987244e-08, 0,
  0, 0, 2.987244e-08, 0.0001530009, 0.000663551, 0.0009392853, 0.000663551, 
    0.0001530009, 2.987244e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 2.636911e-13, 2.989526e-08, 0.0001574448, 0.0006880676, 0.0009750733, 
    0.0006880676, 0.0001574448, 2.989526e-08, 2.636911e-13, 0,
  0, 2.989526e-08, 0.000526949, 0.1337101, 0.206512, 0.2254292, 0.206512, 
    0.1337101, 0.000526949, 2.989526e-08, 0,
  0, 0.0001574448, 0.1337101, 0.2421545, 0.2876507, 0.3013995, 0.2876507, 
    0.2421545, 0.1337101, 0.0001574448, 0,
  0, 0.0006880676, 0.206512, 0.2876507, 0.3281707, 0.3410146, 0.3281707, 
    0.2876507, 0.206512, 0.0006880676, 0,
  0, 0.0009750733, 0.2254292, 0.3013995, 0.3410146, 0.3534367, 0.3410146, 
    0.3013995, 0.2254292, 0.0009750733, 0,
  0, 0.0006880676, 0.206512, 0.2876507, 0.3281707, 0.3410146, 0.3281707, 
    0.2876507, 0.206512, 0.0006880676, 0,
  0, 0.0001574448, 0.1337101, 0.2421545, 0.2876507, 0.3013995, 0.2876507, 
    0.2421545, 0.1337101, 0.0001574448, 0,
  0, 2.989526e-08, 0.000526949, 0.1337101, 0.206512, 0.2254292, 0.206512, 
    0.1337101, 0.000526949, 2.989526e-08, 0,
  0, 2.636912e-13, 2.989527e-08, 0.0001574449, 0.0006880677, 0.0009750734, 
    0.0006880675, 0.0001574447, 2.989528e-08, 2.63691e-13, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 usurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.1325216, 0.2058042, 0.2249885, 0.2058042, 0.1325216, 0, 0, 0,
  0, 0, 0.1325216, 0.2426609, 0.289271, 0.3032196, 0.289271, 0.2426609, 
    0.1325216, 0, 0,
  0, 0, 0.2058042, 0.289271, 0.3293495, 0.3416658, 0.3293495, 0.289271, 
    0.2058042, 0, 0,
  0, 0, 0.2249885, 0.3032196, 0.3416658, 0.3535534, 0.3416658, 0.3032196, 
    0.2249885, 0, 0,
  0, 0, 0.2058042, 0.289271, 0.3293495, 0.3416658, 0.3293495, 0.289271, 
    0.2058042, 0, 0,
  0, 0, 0.1325216, 0.2426609, 0.289271, 0.3032196, 0.289271, 0.2426609, 
    0.1325216, 0, 0,
  0, 0, 0, 0.1325216, 0.2058042, 0.2249885, 0.2058042, 0.1325216, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 3.201627e-05, 0.0002929367, 0.0005178058, 0.0002929367, 
    3.201627e-05, 0, 0, 0,
  0, 0, 5.686403e-05, 0.1326432, 0.2056712, 0.2245772, 0.2056712, 0.1326432, 
    5.686403e-05, 0, 0,
  0, 3.201627e-05, 0.1326432, 0.242601, 0.2890971, 0.3030184, 0.2890971, 
    0.242601, 0.1326432, 3.201627e-05, 0,
  0, 0.0002929367, 0.2056712, 0.2890971, 0.3292324, 0.3416044, 0.3292324, 
    0.2890971, 0.2056712, 0.0002929367, 0,
  0, 0.0005178058, 0.2245772, 0.3030184, 0.3416044, 0.3535409, 0.3416044, 
    0.3030184, 0.2245772, 0.0005178058, 0,
  0, 0.0002929367, 0.2056712, 0.2890971, 0.3292324, 0.3416044, 0.3292324, 
    0.2890971, 0.2056712, 0.0002929367, 0,
  0, 3.201627e-05, 0.1326432, 0.242601, 0.2890971, 0.3030184, 0.2890971, 
    0.242601, 0.1326432, 3.201627e-05, 0,
  0, 0, 5.686403e-05, 0.1326432, 0.2056712, 0.2245772, 0.2056712, 0.1326432, 
    5.686403e-05, 0, 0,
  0, 0, 0, 3.201627e-05, 0.0002929367, 0.0005178058, 0.0002929367, 
    3.201627e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3.499507e-10, 6.994776e-05, 0.0004022547, 0.0006260089, 0.0004022547, 
    6.994776e-05, 3.499507e-10, 0, 0,
  0, 3.499507e-10, 0.0001142617, 0.1327566, 0.205702, 0.2246232, 0.205702, 
    0.1327566, 0.0001142617, 3.499507e-10, 0,
  0, 6.994776e-05, 0.1327566, 0.2425436, 0.2889217, 0.302815, 0.2889217, 
    0.2425436, 0.1327566, 6.994776e-05, 0,
  0, 0.0004022547, 0.205702, 0.2889217, 0.3291154, 0.3415415, 0.3291154, 
    0.2889217, 0.205702, 0.0004022547, 0,
  0, 0.0006260089, 0.2246232, 0.302815, 0.3415415, 0.3535296, 0.3415415, 
    0.302815, 0.2246232, 0.0006260089, 0,
  0, 0.0004022547, 0.205702, 0.2889217, 0.3291154, 0.3415415, 0.3291154, 
    0.2889217, 0.205702, 0.0004022547, 0,
  0, 6.994776e-05, 0.1327566, 0.2425436, 0.2889217, 0.302815, 0.2889217, 
    0.2425436, 0.1327566, 6.994776e-05, 0,
  0, 3.499507e-10, 0.0001142617, 0.1327566, 0.205702, 0.2246232, 0.205702, 
    0.1327566, 0.0001142617, 3.499507e-10, 0,
  0, 0, 3.499507e-10, 6.994776e-05, 0.0004022547, 0.0006260089, 0.0004022547, 
    6.994776e-05, 3.499507e-10, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.146815e-09, 0.0001080381, 0.0005117886, 0.0007343993, 0.0005117886, 
    0.0001080381, 1.146815e-09, 0, 0,
  0, 1.146815e-09, 0.0001718189, 0.1328695, 0.2057316, 0.224668, 0.2057316, 
    0.1328695, 0.0001718189, 1.146815e-09, 0,
  0, 0.0001080381, 0.1328695, 0.2424858, 0.2887474, 0.3026132, 0.2887474, 
    0.2424858, 0.1328695, 0.0001080381, 0,
  0, 0.0005117886, 0.2057316, 0.2887474, 0.3289987, 0.3414782, 0.3289987, 
    0.2887474, 0.2057316, 0.0005117886, 0,
  0, 0.0007343993, 0.224668, 0.3026132, 0.3414782, 0.3535181, 0.3414782, 
    0.3026132, 0.224668, 0.0007343993, 0,
  0, 0.0005117886, 0.2057316, 0.2887474, 0.3289987, 0.3414782, 0.3289987, 
    0.2887474, 0.2057316, 0.0005117886, 0,
  0, 0.0001080381, 0.1328695, 0.2424858, 0.2887474, 0.3026132, 0.2887474, 
    0.2424858, 0.1328695, 0.0001080381, 0,
  0, 1.146815e-09, 0.0001718189, 0.1328695, 0.2057316, 0.224668, 0.2057316, 
    0.1328695, 0.0001718189, 1.146815e-09, 0,
  0, 0, 1.146815e-09, 0.0001080381, 0.0005117886, 0.0007343993, 0.0005117886, 
    0.0001080381, 1.146815e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3.71059e-09, 0.0001152924, 0.0005366366, 0.0007680521, 0.0005366366, 
    0.0001152924, 3.71059e-09, 0, 0,
  0, 3.71059e-09, 0.0002283403, 0.1329929, 0.2058461, 0.2247803, 0.2058461, 
    0.1329929, 0.0002283403, 3.71059e-09, 0,
  0, 0.0001152924, 0.1329929, 0.2424286, 0.2885876, 0.3024359, 0.2885876, 
    0.2424286, 0.1329929, 0.0001152924, 0,
  0, 0.0005366366, 0.2058461, 0.2885876, 0.3288787, 0.3414127, 0.3288787, 
    0.2885876, 0.2058461, 0.0005366366, 0,
  0, 0.0007680521, 0.2247803, 0.3024359, 0.3414127, 0.353507, 0.3414127, 
    0.3024359, 0.2247803, 0.0007680521, 0,
  0, 0.0005366366, 0.2058461, 0.2885876, 0.3288787, 0.3414127, 0.3288787, 
    0.2885876, 0.2058461, 0.0005366366, 0,
  0, 0.0001152924, 0.1329929, 0.2424286, 0.2885876, 0.3024359, 0.2885876, 
    0.2424286, 0.1329929, 0.0001152924, 0,
  0, 3.71059e-09, 0.0002283403, 0.1329929, 0.2058461, 0.2247803, 0.2058461, 
    0.1329929, 0.0002283403, 3.71059e-09, 0,
  0, 0, 3.71059e-09, 0.0001152924, 0.0005366366, 0.0007680521, 0.0005366366, 
    0.0001152924, 3.71059e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 7.089051e-09, 0.000122646, 0.0005616767, 0.0008019177, 0.0005616767, 
    0.000122646, 7.089051e-09, 0, 0,
  0, 7.089051e-09, 0.0002850269, 0.1331159, 0.2059595, 0.2248914, 0.2059595, 
    0.1331159, 0.0002850269, 7.089051e-09, 0,
  0, 0.000122646, 0.1331159, 0.2423711, 0.2884287, 0.30226, 0.2884287, 
    0.2423711, 0.1331159, 0.000122646, 0,
  0, 0.0005616767, 0.2059595, 0.2884287, 0.328759, 0.3413469, 0.328759, 
    0.2884287, 0.2059595, 0.0005616767, 0,
  0, 0.0008019177, 0.2248914, 0.30226, 0.3413469, 0.3534958, 0.3413469, 
    0.30226, 0.2248914, 0.0008019177, 0,
  0, 0.0005616767, 0.2059595, 0.2884287, 0.328759, 0.3413469, 0.328759, 
    0.2884287, 0.2059595, 0.0005616767, 0,
  0, 0.000122646, 0.1331159, 0.2423711, 0.2884287, 0.30226, 0.2884287, 
    0.2423711, 0.1331159, 0.000122646, 0,
  0, 7.089051e-09, 0.0002850269, 0.1331159, 0.2059595, 0.2248914, 0.2059595, 
    0.1331159, 0.0002850269, 7.089051e-09, 0,
  0, 0, 7.089051e-09, 0.000122646, 0.0005616767, 0.0008019177, 0.0005616767, 
    0.000122646, 7.089051e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.134039e-08, 0.0001300937, 0.0005868892, 0.0008359754, 0.0005868892, 
    0.0001300937, 1.134039e-08, 0, 0,
  0, 1.134039e-08, 0.0003418765, 0.1332385, 0.206072, 0.2250013, 0.206072, 
    0.1332385, 0.0003418765, 1.134039e-08, 0,
  0, 0.0001300937, 0.1332385, 0.2423133, 0.2882708, 0.3020855, 0.2882708, 
    0.2423133, 0.1332385, 0.0001300937, 0,
  0, 0.0005868892, 0.206072, 0.2882708, 0.3286397, 0.3412811, 0.3286397, 
    0.2882708, 0.206072, 0.0005868892, 0,
  0, 0.0008359754, 0.2250013, 0.3020855, 0.3412811, 0.3534843, 0.3412811, 
    0.3020855, 0.2250013, 0.0008359754, 0,
  0, 0.0005868892, 0.206072, 0.2882708, 0.3286397, 0.3412811, 0.3286397, 
    0.2882708, 0.206072, 0.0005868892, 0,
  0, 0.0001300937, 0.1332385, 0.2423133, 0.2882708, 0.3020855, 0.2882708, 
    0.2423133, 0.1332385, 0.0001300937, 0,
  0, 1.134039e-08, 0.0003418765, 0.1332385, 0.206072, 0.2250013, 0.206072, 
    0.1332385, 0.0003418765, 1.134039e-08, 0,
  0, 0, 1.134039e-08, 0.0001300937, 0.0005868892, 0.0008359754, 0.0005868892, 
    0.0001300937, 1.134039e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.651755e-08, 0.0001376354, 0.0006122729, 0.0008702234, 0.0006122729, 
    0.0001376354, 1.651755e-08, 0, 0,
  0, 1.651755e-08, 0.0003988868, 0.1333608, 0.2061835, 0.22511, 0.2061835, 
    0.1333608, 0.0003988868, 1.651755e-08, 0,
  0, 0.0001376354, 0.1333608, 0.2422552, 0.2881137, 0.3019123, 0.2881137, 
    0.2422552, 0.1333608, 0.0001376354, 0,
  0, 0.0006122729, 0.2061835, 0.2881137, 0.3285207, 0.341215, 0.3285207, 
    0.2881137, 0.2061835, 0.0006122729, 0,
  0, 0.0008702234, 0.22511, 0.3019123, 0.341215, 0.3534726, 0.341215, 
    0.3019123, 0.22511, 0.0008702234, 0,
  0, 0.0006122729, 0.2061835, 0.2881137, 0.3285207, 0.341215, 0.3285207, 
    0.2881137, 0.2061835, 0.0006122729, 0,
  0, 0.0001376354, 0.1333608, 0.2422552, 0.2881137, 0.3019123, 0.2881137, 
    0.2422552, 0.1333608, 0.0001376354, 0,
  0, 1.651755e-08, 0.0003988868, 0.1333608, 0.2061835, 0.22511, 0.2061835, 
    0.1333608, 0.0003988868, 1.651755e-08, 0,
  0, 0, 1.651755e-08, 0.0001376354, 0.0006122729, 0.0008702234, 0.0006122729, 
    0.0001376354, 1.651755e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 2.267689e-08, 0.0001452712, 0.0006378272, 0.0009046606, 0.0006378272, 
    0.0001452712, 2.267689e-08, 0, 0,
  0, 2.267689e-08, 0.0004560562, 0.1334826, 0.206294, 0.2252176, 0.206294, 
    0.1334826, 0.0004560562, 2.267689e-08, 0,
  0, 0.0001452712, 0.1334826, 0.2421968, 0.2879576, 0.3017404, 0.2879576, 
    0.2421968, 0.1334826, 0.0001452712, 0,
  0, 0.0006378272, 0.206294, 0.2879576, 0.3284021, 0.3411488, 0.3284021, 
    0.2879576, 0.206294, 0.0006378272, 0,
  0, 0.0009046606, 0.2252176, 0.3017404, 0.3411488, 0.3534607, 0.3411488, 
    0.3017404, 0.2252176, 0.0009046606, 0,
  0, 0.0006378272, 0.206294, 0.2879576, 0.3284021, 0.3411488, 0.3284021, 
    0.2879576, 0.206294, 0.0006378272, 0,
  0, 0.0001452712, 0.1334826, 0.2421968, 0.2879576, 0.3017404, 0.2879576, 
    0.2421968, 0.1334826, 0.0001452712, 0,
  0, 2.267689e-08, 0.0004560562, 0.1334826, 0.206294, 0.2252176, 0.206294, 
    0.1334826, 0.0004560562, 2.267689e-08, 0,
  0, 0, 2.267689e-08, 0.0001452712, 0.0006378272, 0.0009046606, 0.0006378272, 
    0.0001452712, 2.267689e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 2.987244e-08, 0.0001530009, 0.000663551, 0.0009392853, 0.000663551, 
    0.0001530009, 2.987244e-08, 0, 0,
  0, 2.987244e-08, 0.0005133827, 0.1336041, 0.2064035, 0.2253239, 0.2064035, 
    0.1336041, 0.0005133827, 2.987244e-08, 0,
  0, 0.0001530009, 0.1336041, 0.2421382, 0.2878024, 0.3015697, 0.2878024, 
    0.2421382, 0.1336041, 0.0001530009, 0,
  0, 0.000663551, 0.2064035, 0.2878024, 0.3282839, 0.3410824, 0.3282839, 
    0.2878024, 0.2064035, 0.000663551, 0,
  0, 0.0009392853, 0.2253239, 0.3015697, 0.3410824, 0.3534486, 0.3410824, 
    0.3015697, 0.2253239, 0.0009392853, 0,
  0, 0.000663551, 0.2064035, 0.2878024, 0.3282839, 0.3410824, 0.3282839, 
    0.2878024, 0.2064035, 0.000663551, 0,
  0, 0.0001530009, 0.1336041, 0.2421382, 0.2878024, 0.3015697, 0.2878024, 
    0.2421382, 0.1336041, 0.0001530009, 0,
  0, 2.987244e-08, 0.0005133827, 0.1336041, 0.2064035, 0.2253239, 0.2064035, 
    0.1336041, 0.0005133827, 2.987244e-08, 0,
  0, 0, 2.987244e-08, 0.0001530009, 0.000663551, 0.0009392853, 0.000663551, 
    0.0001530009, 2.987244e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 2.636911e-13, 2.989526e-08, 0.0001574448, 0.0006880676, 0.0009750733, 
    0.0006880676, 0.0001574448, 2.989526e-08, 2.636911e-13, 0,
  0, 2.989526e-08, 0.000526949, 0.1337101, 0.206512, 0.2254292, 0.206512, 
    0.1337101, 0.000526949, 2.989526e-08, 0,
  0, 0.0001574448, 0.1337101, 0.2421545, 0.2876507, 0.3013995, 0.2876507, 
    0.2421545, 0.1337101, 0.0001574448, 0,
  0, 0.0006880676, 0.206512, 0.2876507, 0.3281707, 0.3410146, 0.3281707, 
    0.2876507, 0.206512, 0.0006880676, 0,
  0, 0.0009750733, 0.2254292, 0.3013995, 0.3410146, 0.3534367, 0.3410146, 
    0.3013995, 0.2254292, 0.0009750733, 0,
  0, 0.0006880676, 0.206512, 0.2876507, 0.3281707, 0.3410146, 0.3281707, 
    0.2876507, 0.206512, 0.0006880676, 0,
  0, 0.0001574448, 0.1337101, 0.2421545, 0.2876507, 0.3013995, 0.2876507, 
    0.2421545, 0.1337101, 0.0001574448, 0,
  0, 2.989526e-08, 0.000526949, 0.1337101, 0.206512, 0.2254292, 0.206512, 
    0.1337101, 0.000526949, 2.989526e-08, 0,
  0, 2.636911e-13, 2.989526e-08, 0.0001574448, 0.0006880676, 0.0009750733, 
    0.0006880676, 0.0001574448, 2.989526e-08, 2.636911e-13, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 uvel =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -0.0003132102, -0.003165813, -0.003779339, 0.003779339, 0.003165813, 
    0.0003132102, 0, 0,
  0, 0.0008256877, -0.008360734, -0.005990916, -0.002186223, 0.002186223, 
    0.005990916, 0.008360734, -0.0008256877, 0,
  0, -0.01155192, -0.00988832, -0.004564836, -0.0007603604, 0.0007603604, 
    0.004564836, 0.00988832, 0.01155192, 0,
  0, -0.0525986, -0.01105339, -0.002173914, -0.0001664206, 0.0001664206, 
    0.002173914, 0.01105339, 0.0525986, 0,
  0, -0.0525986, -0.01105339, -0.002173914, -0.0001664206, 0.0001664206, 
    0.002173914, 0.01105339, 0.0525986, 0,
  0, -0.01155192, -0.00988832, -0.004564836, -0.0007603604, 0.0007603604, 
    0.004564836, 0.00988832, 0.01155192, 0,
  0, 0.0008256877, -0.008360734, -0.005990916, -0.002186223, 0.002186223, 
    0.005990916, 0.008360734, -0.0008256877, 0,
  0, 0, -0.0003132102, -0.003165813, -0.003779339, 0.003779339, 0.003165813, 
    0.0003132102, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -0.000247678, -0.003127966, -0.003727764, 0.003727764, 0.003127966, 
    0.000247678, 0, 0,
  0, 0.0008988078, -0.008286852, -0.005943459, -0.002137286, 0.002137286, 
    0.005943459, 0.008286852, -0.0008988078, 0,
  0, -0.01142125, -0.009812617, -0.004470771, -0.000737313, 0.000737313, 
    0.004470771, 0.009812617, 0.01142125, 0,
  0, -0.05188848, -0.01079278, -0.002120323, -0.0001542805, 0.0001542805, 
    0.002120323, 0.01079278, 0.05188848, 0,
  0, -0.05188848, -0.01079278, -0.002120323, -0.0001542805, 0.0001542805, 
    0.002120323, 0.01079278, 0.05188848, 0,
  0, -0.01142125, -0.009812617, -0.004470771, -0.000737313, 0.000737313, 
    0.004470771, 0.009812617, 0.01142125, 0,
  0, 0.0008988078, -0.008286852, -0.005943459, -0.002137286, 0.002137286, 
    0.005943459, 0.008286852, -0.0008988078, 0,
  0, 0, -0.000247678, -0.003127966, -0.003727764, 0.003727764, 0.003127966, 
    0.000247678, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -0.0001338964, -0.003009181, -0.00357941, 0.00357941, 0.003009181, 
    0.0001338964, 0, 0,
  0, 0.001005922, -0.008015784, -0.005748612, -0.001999517, 0.001999517, 
    0.005748612, 0.008015784, -0.001005922, 0,
  0, -0.01098942, -0.00950125, -0.004218965, -0.000681401, 0.000681401, 
    0.004218965, 0.00950125, 0.01098942, 0,
  0, -0.04981515, -0.01007572, -0.001982236, -0.0001292175, 0.0001292175, 
    0.001982236, 0.01007572, 0.04981515, 0,
  0, -0.04981515, -0.01007572, -0.001982236, -0.0001292175, 0.0001292175, 
    0.001982236, 0.01007572, 0.04981515, 0,
  0, -0.01098942, -0.00950125, -0.004218965, -0.000681401, 0.000681401, 
    0.004218965, 0.00950125, 0.01098942, 0,
  0, 0.001005922, -0.008015784, -0.005748612, -0.001999517, 0.001999517, 
    0.005748612, 0.008015784, -0.001005922, 0,
  0, 0, -0.0001338964, -0.003009181, -0.00357941, 0.00357941, 0.003009181, 
    0.0001338964, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -4.092442e-05, -0.002763917, -0.003310581, 0.003310581, 0.002763917, 
    4.092442e-05, 0, 0,
  0, 0.001032454, -0.007404672, -0.005318087, -0.001799537, 0.001799537, 
    0.005318087, 0.007404672, -0.001032454, 0,
  0, -0.01008927, -0.00879538, -0.003830721, -0.0006064072, 0.0006064072, 
    0.003830721, 0.00879538, 0.01008927, 0,
  0, -0.04598061, -0.009030757, -0.001783949, -0.0001023342, 0.0001023342, 
    0.001783949, 0.009030757, 0.04598061, 0,
  0, -0.04598061, -0.009030757, -0.001783949, -0.0001023342, 0.0001023342, 
    0.001783949, 0.009030757, 0.04598061, 0,
  0, -0.01008927, -0.00879538, -0.003830721, -0.0006064072, 0.0006064072, 
    0.003830721, 0.00879538, 0.01008927, 0,
  0, 0.001032454, -0.007404672, -0.005318087, -0.001799537, 0.001799537, 
    0.005318087, 0.007404672, -0.001032454, 0,
  0, 0, -4.092442e-05, -0.002763917, -0.003310581, 0.003310581, 0.002763917, 
    4.092442e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.882779e-05, -0.002400004, -0.002906606, 0.002906606, 0.002400004, 
    -1.882779e-05, 0, 0,
  0, 0.0009651849, -0.006466162, -0.004651948, -0.001546011, 0.001546011, 
    0.004651948, 0.006466162, -0.0009651849, 0,
  0, -0.008752258, -0.007693929, -0.003310903, -0.0005176318, 0.0005176318, 
    0.003310903, 0.007693929, 0.008752258, 0,
  0, -0.04026955, -0.00771859, -0.001535694, -7.849183e-05, 7.849183e-05, 
    0.001535694, 0.00771859, 0.04026955, 0,
  0, -0.04026955, -0.00771859, -0.001535694, -7.849183e-05, 7.849183e-05, 
    0.001535694, 0.00771859, 0.04026955, 0,
  0, -0.008752258, -0.007693929, -0.003310903, -0.0005176318, 0.0005176318, 
    0.003310903, 0.007693929, 0.008752258, 0,
  0, 0.0009651849, -0.006466162, -0.004651948, -0.001546011, 0.001546011, 
    0.004651948, 0.006466162, -0.0009651849, 0,
  0, 0, 1.882779e-05, -0.002400004, -0.002906606, 0.002906606, 0.002400004, 
    -1.882779e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 5.001188e-05, -0.001955896, -0.002395972, 0.002395972, 0.001955896, 
    -5.001188e-05, 0, 0,
  0, 0.0008288237, -0.005296842, -0.003816402, -0.001252671, 0.001252671, 
    0.003816402, 0.005296842, -0.0008288237, 0,
  0, -0.007124439, -0.006310518, -0.002694009, -0.0004183753, 0.0004183753, 
    0.002694009, 0.006310518, 0.007124439, 0,
  0, -0.03311698, -0.006221511, -0.001249252, -5.834021e-05, 5.834021e-05, 
    0.001249252, 0.006221511, 0.03311698, 0,
  0, -0.03311698, -0.006221511, -0.001249252, -5.834021e-05, 5.834021e-05, 
    0.001249252, 0.006221511, 0.03311698, 0,
  0, -0.007124439, -0.006310518, -0.002694009, -0.0004183753, 0.0004183753, 
    0.002694009, 0.006310518, 0.007124439, 0,
  0, 0.0008288237, -0.005296842, -0.003816402, -0.001252671, 0.001252671, 
    0.003816402, 0.005296842, -0.0008288237, 0,
  0, 0, 5.001188e-05, -0.001955896, -0.002395972, 0.002395972, 0.001955896, 
    -5.001188e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 5.845296e-05, -0.001469448, -0.001819022, 0.001819022, 0.001469448, 
    -5.845296e-05, 0, 0,
  0, 0.0006475092, -0.003997323, -0.002883687, -0.0009378714, 0.0009378714, 
    0.002883687, 0.003997323, -0.0006475092, 0,
  0, -0.00534637, -0.004766757, -0.002023412, -0.0003130873, 0.0003130873, 
    0.002023412, 0.004766757, 0.00534637, 0,
  0, -0.02509051, -0.004635514, -0.000939752, -4.102458e-05, 4.102458e-05, 
    0.000939752, 0.004635514, 0.02509051, 0,
  0, -0.02509051, -0.004635514, -0.000939752, -4.102458e-05, 4.102458e-05, 
    0.000939752, 0.004635514, 0.02509051, 0,
  0, -0.00534637, -0.004766757, -0.002023412, -0.0003130873, 0.0003130873, 
    0.002023412, 0.004766757, 0.00534637, 0,
  0, 0.0006475092, -0.003997323, -0.002883687, -0.0009378714, 0.0009378714, 
    0.002883687, 0.003997323, -0.0006475092, 0,
  0, 0, 5.845296e-05, -0.001469448, -0.001819022, 0.001819022, 0.001469448, 
    -5.845296e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 4.978968e-05, -0.0009694969, -0.001211213, 0.001211213, 0.0009694969, 
    -4.978968e-05, 0, 0,
  0, 0.0004403218, -0.002647395, -0.001911809, -0.0006173779, 0.0006173779, 
    0.001911809, 0.002647395, -0.0004403218, 0,
  0, -0.003523594, -0.003159238, -0.00133532, -0.0002061807, 0.0002061807, 
    0.00133532, 0.003159238, 0.003523594, 0,
  0, -0.01667722, -0.003038258, -0.0006215644, -2.578999e-05, 2.578999e-05, 
    0.0006215644, 0.003038258, 0.01667722, 0,
  0, -0.01667722, -0.003038258, -0.0006215644, -2.578999e-05, 2.578999e-05, 
    0.0006215644, 0.003038258, 0.01667722, 0,
  0, -0.003523594, -0.003159238, -0.00133532, -0.0002061807, 0.0002061807, 
    0.00133532, 0.003159238, 0.003523594, 0,
  0, 0.0004403218, -0.002647395, -0.001911809, -0.0006173779, 0.0006173779, 
    0.001911809, 0.002647395, -0.0004403218, 0,
  0, 0, 4.978968e-05, -0.0009694969, -0.001211213, 0.001211213, 0.0009694969, 
    -4.978968e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 2.896606e-05, -0.0004756116, -0.0005989244, 0.0005989244, 
    0.0004756116, -2.896606e-05, 0, 0,
  0, 0.0002212498, -0.001302959, -0.0009417262, -0.0003023877, 0.0003023877, 
    0.0009417262, 0.001302959, -0.0002212498, 0,
  0, -0.001726917, -0.001555736, -0.000655379, -0.0001010627, 0.0001010627, 
    0.000655379, 0.001555736, 0.001726917, 0,
  0, -0.008234199, -0.001482464, -0.0003057959, -1.220087e-05, 1.220087e-05, 
    0.0003057959, 0.001482464, 0.008234199, 0,
  0, -0.008234199, -0.001482464, -0.0003057959, -1.220087e-05, 1.220087e-05, 
    0.0003057959, 0.001482464, 0.008234199, 0,
  0, -0.001726917, -0.001555736, -0.000655379, -0.0001010627, 0.0001010627, 
    0.000655379, 0.001555736, 0.001726917, 0,
  0, 0.0002212498, -0.001302959, -0.0009417262, -0.0003023877, 0.0003023877, 
    0.0009417262, 0.001302959, -0.0002212498, 0,
  0, 0, 2.896606e-05, -0.0004756116, -0.0005989244, 0.0005989244, 
    0.0004756116, -2.896606e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -1.242242e-08, -7.061802e-09, -2.447388e-09, 2.447388e-09, 
    7.061802e-09, 1.242242e-08, 0, 0,
  0, -1.179029e-08, -2.355311e-08, -1.515827e-08, -4.68496e-09, 4.68496e-09, 
    1.515827e-08, 2.355311e-08, 1.179029e-08, 0,
  0, -3.384802e-08, -2.524052e-08, -1.557322e-08, -5.164675e-09, 
    5.164675e-09, 1.557322e-08, 2.524052e-08, 3.384802e-08, 0,
  0, -5.10667e-08, -2.730837e-08, -1.478742e-08, -5.859598e-09, 5.859598e-09, 
    1.478742e-08, 2.730837e-08, 5.10667e-08, 0,
  0, -5.10667e-08, -2.730837e-08, -1.478742e-08, -5.859598e-09, 5.859598e-09, 
    1.478742e-08, 2.730837e-08, 5.10667e-08, 0,
  0, -3.384802e-08, -2.524052e-08, -1.557322e-08, -5.164675e-09, 
    5.164675e-09, 1.557322e-08, 2.524052e-08, 3.384802e-08, 0,
  0, -1.179029e-08, -2.355311e-08, -1.515827e-08, -4.68496e-09, 4.68496e-09, 
    1.515827e-08, 2.355311e-08, 1.179029e-08, 0,
  0, 0, -1.242242e-08, -7.061802e-09, -2.447388e-09, 2.447388e-09, 
    7.061802e-09, 1.242242e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0001409117, -0.0001409117, 0, 0, 0, 0,
  0, 0, -0.0004603508, -0.002767604, -0.0005696231, 0.0005696231, 
    0.002767604, 0.0004603508, 0, 0,
  0, 0.001588732, -0.008342631, -0.006091888, -0.002037874, 0.002037874, 
    0.006091888, 0.008342631, -0.001588732, 0,
  0, -0.01383611, -0.00982201, -0.004516106, -0.0008045277, 0.0008045277, 
    0.004516106, 0.00982201, 0.01383611, 0,
  0.002904966, -0.01093761, -0.01079595, -0.002305073, -0.0001358764, 
    0.0001358764, 0.002305073, 0.01079595, 0.01093761, -0.002904966,
  0.002904966, -0.01093761, -0.01079595, -0.002305073, -0.0001358764, 
    0.0001358764, 0.002305073, 0.01079595, 0.01093761, -0.002904966,
  0, -0.01383611, -0.00982201, -0.004516106, -0.0008045277, 0.0008045277, 
    0.004516106, 0.00982201, 0.01383611, 0,
  0, 0.001588732, -0.008342631, -0.006091888, -0.002037874, 0.002037874, 
    0.006091888, 0.008342631, -0.001588732, 0,
  0, 0, -0.0004603508, -0.002767604, -0.0005696231, 0.0005696231, 
    0.002767604, 0.0004603508, 0, 0,
  0, 0, 0, 0, 0.0001409117, -0.0001409117, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0001418827, -0.0001418827, 0, 0, 0, 0,
  0, 0, -0.0003771874, -0.002750773, -0.0005671459, 0.0005671459, 
    0.002750773, 0.0003771874, 0, 0,
  0, 0.001689613, -0.008274466, -0.006040138, -0.002014322, 0.002014322, 
    0.006040138, 0.008274466, -0.001689613, 0,
  0, -0.01374504, -0.009729467, -0.004426829, -0.0007758784, 0.0007758784, 
    0.004426829, 0.009729467, 0.01374504, 0,
  0.002900456, -0.01086727, -0.01069149, -0.002220682, -0.0001304481, 
    0.0001304481, 0.002220682, 0.01069149, 0.01086727, -0.002900456,
  0.002900456, -0.01086727, -0.01069149, -0.002220682, -0.0001304481, 
    0.0001304481, 0.002220682, 0.01069149, 0.01086727, -0.002900456,
  0, -0.01374504, -0.009729467, -0.004426829, -0.0007758784, 0.0007758784, 
    0.004426829, 0.009729467, 0.01374504, 0,
  0, 0.001689613, -0.008274466, -0.006040138, -0.002014322, 0.002014322, 
    0.006040138, 0.008274466, -0.001689613, 0,
  0, 0, -0.0003771874, -0.002750773, -0.0005671459, 0.0005671459, 
    0.002750773, 0.0003771874, 0, 0,
  0, 0, 0, 0, 0.0001418827, -0.0001418827, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0001375639, -0.0001375639, 0, 0, 0, 0,
  0, 0, -0.0002335275, -0.00267804, -0.0005429088, 0.0005429088, 0.00267804, 
    0.0002335275, 0, 0,
  0, 0.001813428, -0.008012175, -0.005836438, -0.001930867, 0.001930867, 
    0.005836438, 0.008012175, -0.001813428, 0,
  0, -0.01332963, -0.009390969, -0.004183661, -0.0007077734, 0.0007077734, 
    0.004183661, 0.009390969, 0.01332963, 0,
  0.002809787, -0.01050294, -0.01026892, -0.002026674, -0.000116664, 
    0.000116664, 0.002026674, 0.01026892, 0.01050294, -0.002809787,
  0.002809787, -0.01050294, -0.01026892, -0.002026674, -0.000116664, 
    0.000116664, 0.002026674, 0.01026892, 0.01050294, -0.002809787,
  0, -0.01332963, -0.009390969, -0.004183661, -0.0007077734, 0.0007077734, 
    0.004183661, 0.009390969, 0.01332963, 0,
  0, 0.001813428, -0.008012175, -0.005836438, -0.001930867, 0.001930867, 
    0.005836438, 0.008012175, -0.001813428, 0,
  0, 0, -0.0002335275, -0.00267804, -0.0005429088, 0.0005429088, 0.00267804, 
    0.0002335275, 0, 0,
  0, 0, 0, 0, 0.0001375639, -0.0001375639, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0001255195, -0.0001255195, 0, 0, 0, 0,
  0, 0, -0.0001143945, -0.002484142, -0.00049014, 0.00049014, 0.002484142, 
    0.0001143945, 0, 0,
  0, 0.001808339, -0.007412508, -0.005389567, -0.001774436, 0.001774436, 
    0.005389567, 0.007412508, -0.001808339, 0,
  0, -0.01232277, -0.008663377, -0.003806251, -0.0006214951, 0.0006214951, 
    0.003806251, 0.008663377, 0.01232277, 0,
  0.002591708, -0.009678153, -0.009446746, -0.001783908, -9.855127e-05, 
    9.855127e-05, 0.001783908, 0.009446746, 0.009678153, -0.002591708,
  0.002591708, -0.009678153, -0.009446746, -0.001783908, -9.855127e-05, 
    9.855127e-05, 0.001783908, 0.009446746, 0.009678153, -0.002591708,
  0, -0.01232277, -0.008663377, -0.003806251, -0.0006214951, 0.0006214951, 
    0.003806251, 0.008663377, 0.01232277, 0,
  0, 0.001808339, -0.007412508, -0.005389567, -0.001774436, 0.001774436, 
    0.005389567, 0.007412508, -0.001808339, 0,
  0, 0, -0.0001143945, -0.002484142, -0.00049014, 0.00049014, 0.002484142, 
    0.0001143945, 0, 0,
  0, 0, 0, 0, 0.0001255195, -0.0001255195, 0, 0, 0, 0,
  0, 0, 0, 0, 0.000107753, -0.000107753, 0, 0, 0, 0,
  0, 0, -3.382427e-05, -0.002175087, -0.0004169835, 0.0004169835, 
    0.002175087, 3.382427e-05, 0, 0,
  0, 0.001664641, -0.006482529, -0.004706029, -0.001546509, 0.001546509, 
    0.004706029, 0.006482529, -0.001664641, 0,
  0, -0.01076163, -0.007557421, -0.003295617, -0.0005249813, 0.0005249813, 
    0.003295617, 0.007557421, 0.01076163, 0,
  0.002257105, -0.008424691, -0.008239493, -0.001509017, -7.993602e-05, 
    7.993602e-05, 0.001509017, 0.008239493, 0.008424691, -0.002257105,
  0.002257105, -0.008424691, -0.008239493, -0.001509017, -7.993602e-05, 
    7.993602e-05, 0.001509017, 0.008239493, 0.008424691, -0.002257105,
  0, -0.01076163, -0.007557421, -0.003295617, -0.0005249813, 0.0005249813, 
    0.003295617, 0.007557421, 0.01076163, 0,
  0, 0.001664641, -0.006482529, -0.004706029, -0.001546509, 0.001546509, 
    0.004706029, 0.006482529, -0.001664641, 0,
  0, 0, -3.382427e-05, -0.002175087, -0.0004169835, 0.0004169835, 
    0.002175087, 3.382427e-05, 0, 0,
  0, 0, 0, 0, 0.000107753, -0.000107753, 0, 0, 0, 0,
  0, 0, 0, 0, 8.679642e-05, -8.679642e-05, 0, 0, 0, 0,
  0, 0, 1.36996e-05, -0.001785389, -0.0003332556, 0.0003332556, 0.001785389, 
    -1.36996e-05, 0, 0,
  0, 0.001416857, -0.005317794, -0.003855044, -0.001266169, 0.001266169, 
    0.003855044, 0.005317794, -0.001416857, 0,
  0, -0.008815134, -0.006185435, -0.0026857, -0.0004209878, 0.0004209878, 
    0.0026857, 0.006185435, 0.008815134, 0,
  0.001843565, -0.006879662, -0.006750421, -0.00121061, -6.231098e-05, 
    6.231098e-05, 0.00121061, 0.006750421, 0.006879662, -0.001843565,
  0.001843565, -0.006879662, -0.006750421, -0.00121061, -6.231098e-05, 
    6.231098e-05, 0.00121061, 0.006750421, 0.006879662, -0.001843565,
  0, -0.008815134, -0.006185435, -0.0026857, -0.0004209878, 0.0004209878, 
    0.0026857, 0.006185435, 0.008815134, 0,
  0, 0.001416857, -0.005317794, -0.003855044, -0.001266169, 0.001266169, 
    0.003855044, 0.005317794, -0.001416857, 0,
  0, 0, 1.36996e-05, -0.001785389, -0.0003332556, 0.0003332556, 0.001785389, 
    -1.36996e-05, 0, 0,
  0, 0, 0, 0, 8.679642e-05, -8.679642e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 6.454564e-05, -6.454564e-05, 0, 0, 0, 0,
  0, 0, 3.488674e-05, -0.001349935, -0.0002460758, 0.0002460758, 0.001349935, 
    -3.488674e-05, 0, 0,
  0, 0.001100926, -0.004019278, -0.0029098, -0.0009557179, 0.0009557179, 
    0.0029098, 0.004019278, -0.001100926, 0,
  0, -0.00665365, -0.004665238, -0.002020023, -0.0003131764, 0.0003131764, 
    0.002020023, 0.004665238, 0.00665365, 0,
  0.00138761, -0.00517776, -0.005098342, -0.0009005336, -4.56211e-05, 
    4.56211e-05, 0.0009005336, 0.005098342, 0.00517776, -0.00138761,
  0.00138761, -0.00517776, -0.005098342, -0.0009005336, -4.56211e-05, 
    4.56211e-05, 0.0009005336, 0.005098342, 0.00517776, -0.00138761,
  0, -0.00665365, -0.004665238, -0.002020023, -0.0003131764, 0.0003131764, 
    0.002020023, 0.004665238, 0.00665365, 0,
  0, 0.001100926, -0.004019278, -0.0029098, -0.0009557179, 0.0009557179, 
    0.0029098, 0.004019278, -0.001100926, 0,
  0, 0, 3.488674e-05, -0.001349935, -0.0002460758, 0.0002460758, 0.001349935, 
    -3.488674e-05, 0, 0,
  0, 0, 0, 0, 6.454564e-05, -6.454564e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 4.223891e-05, -4.223891e-05, 0, 0, 0, 0,
  0, 0, 3.609539e-05, -0.0008961188, -0.0001599589, 0.0001599589, 
    0.0008961188, -3.609539e-05, 0, 0,
  0, 0.0007463105, -0.002667287, -0.001928339, -0.0006334924, 0.0006334924, 
    0.001928339, 0.002667287, -0.0007463105, 0,
  0, -0.004410344, -0.003089655, -0.001335082, -0.0002053431, 0.0002053431, 
    0.001335082, 0.003089655, 0.004410344, 0,
  0.0009171122, -0.003422141, -0.003381234, -0.0005902908, -2.968416e-05, 
    2.968416e-05, 0.0005902908, 0.003381234, 0.003422141, -0.0009171122,
  0.0009171122, -0.003422141, -0.003381234, -0.0005902908, -2.968416e-05, 
    2.968416e-05, 0.0005902908, 0.003381234, 0.003422141, -0.0009171122,
  0, -0.004410344, -0.003089655, -0.001335082, -0.0002053431, 0.0002053431, 
    0.001335082, 0.003089655, 0.004410344, 0,
  0, 0.0007463105, -0.002667287, -0.001928339, -0.0006334924, 0.0006334924, 
    0.001928339, 0.002667287, -0.0007463105, 0,
  0, 0, 3.609539e-05, -0.0008961188, -0.0001599589, 0.0001599589, 
    0.0008961188, -3.609539e-05, 0, 0,
  0, 0, 0, 0, 4.223891e-05, -4.223891e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 2.061441e-05, -2.061441e-05, 0, 0, 0, 0,
  0, 0, 2.297726e-05, -0.0004427537, -7.752377e-05, 7.752377e-05, 
    0.0004427537, -2.297726e-05, 0, 0,
  0, 0.000374839, -0.001317347, -0.0009509482, -0.0003124892, 0.0003124892, 
    0.0009509482, 0.001317347, -0.000374839, 0,
  0, -0.002176257, -0.001522762, -0.000656846, -0.0001004071, 0.0001004071, 
    0.000656846, 0.001522762, 0.002176257, 0,
  0.000450985, -0.001682918, -0.001668764, -0.0002885073, -1.447968e-05, 
    1.447968e-05, 0.0002885073, 0.001668764, 0.001682918, -0.000450985,
  0.000450985, -0.001682918, -0.001668764, -0.0002885073, -1.447968e-05, 
    1.447968e-05, 0.0002885073, 0.001668764, 0.001682918, -0.000450985,
  0, -0.002176257, -0.001522762, -0.000656846, -0.0001004071, 0.0001004071, 
    0.000656846, 0.001522762, 0.002176257, 0,
  0, 0.000374839, -0.001317347, -0.0009509482, -0.0003124892, 0.0003124892, 
    0.0009509482, 0.001317347, -0.000374839, 0,
  0, 0, 2.297726e-05, -0.0004427537, -7.752377e-05, 7.752377e-05, 
    0.0004427537, -2.297726e-05, 0, 0,
  0, 0, 0, 0, 2.061441e-05, -2.061441e-05, 0, 0, 0, 0,
  0, 0, 0, 0, -3.758351e-10, 3.758351e-10, 0, 0, 0, 0,
  0, 0, -1.267312e-08, -6.30858e-09, -2.031621e-09, 2.031621e-09, 
    6.30858e-09, 1.267312e-08, 0, 0,
  0, -1.173665e-08, -2.343477e-08, -1.545185e-08, -4.982604e-09, 
    4.982604e-09, 1.545185e-08, 2.343477e-08, 1.173665e-08, 0,
  0, -3.397699e-08, -2.529044e-08, -1.544368e-08, -5.082978e-09, 
    5.082978e-09, 1.544368e-08, 2.529044e-08, 3.397699e-08, 0,
  8.236872e-09, -3.650524e-08, -2.602708e-08, -1.528052e-08, -5.71314e-09, 
    5.71314e-09, 1.528052e-08, 2.602708e-08, 3.650524e-08, -8.236872e-09,
  8.236872e-09, -3.650524e-08, -2.602708e-08, -1.528052e-08, -5.71314e-09, 
    5.71314e-09, 1.528052e-08, 2.602708e-08, 3.650524e-08, -8.236872e-09,
  0, -3.397699e-08, -2.529044e-08, -1.544368e-08, -5.082978e-09, 
    5.082978e-09, 1.544368e-08, 2.529044e-08, 3.397699e-08, 0,
  0, -1.173665e-08, -2.343477e-08, -1.545185e-08, -4.982604e-09, 
    4.982604e-09, 1.545185e-08, 2.343477e-08, 1.173665e-08, 0,
  0, 0, -1.267312e-08, -6.30858e-09, -2.031621e-09, 2.031621e-09, 
    6.30858e-09, 1.267312e-08, 0, 0,
  0, 0, 0, 0, -3.758351e-10, 3.758351e-10, 0, 0, 0, 0,
  0, 0, 0, 0, 0.000141204, -0.000141204, 0, 0, 0, 0,
  0, 0, -0.0004718868, -0.002775271, -0.0005710098, 0.0005710098, 
    0.002775271, 0.0004718868, 0, 0,
  0, 0.001573083, -0.008346623, -0.006071293, -0.002029181, 0.002029181, 
    0.006071293, 0.008346623, -0.001573083, 0,
  0, -0.01385412, -0.009787603, -0.004500326, -0.0008072912, 0.0008072912, 
    0.004500326, 0.009787603, 0.01385412, 0,
  0.002907086, -0.01094661, -0.01073877, -0.002313738, -0.0001384091, 
    0.0001384091, 0.002313738, 0.01073877, 0.01094661, -0.002907086,
  0.002907086, -0.01094661, -0.01073877, -0.002313738, -0.0001384091, 
    0.0001384091, 0.002313738, 0.01073877, 0.01094661, -0.002907086,
  0, -0.01385412, -0.009787603, -0.004500326, -0.0008072912, 0.0008072912, 
    0.004500326, 0.009787603, 0.01385412, 0,
  0, 0.001573083, -0.008346623, -0.006071293, -0.002029181, 0.002029181, 
    0.006071293, 0.008346623, -0.001573083, 0,
  0, 0, -0.0004718868, -0.002775271, -0.0005710098, 0.0005710098, 
    0.002775271, 0.0004718868, 0, 0,
  0, 0, 0, 0, 0.000141204, -0.000141204, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0001421608, -0.0001421608, 0, 0, 0, 0,
  0, 0, -0.000388854, -0.002758372, -0.0005684611, 0.0005684611, 0.002758372, 
    0.000388854, 0, 0,
  0, 0.001673691, -0.008278607, -0.006019558, -0.00200568, 0.00200568, 
    0.006019558, 0.008278607, -0.001673691, 0,
  0, -0.01376272, -0.00969515, -0.004411527, -0.0007787212, 0.0007787212, 
    0.004411527, 0.00969515, 0.01376272, 0,
  0.002902497, -0.01087582, -0.01063459, -0.002229519, -0.0001328241, 
    0.0001328241, 0.002229519, 0.01063459, 0.01087582, -0.002902497,
  0.002902497, -0.01087582, -0.01063459, -0.002229519, -0.0001328241, 
    0.0001328241, 0.002229519, 0.01063459, 0.01087582, -0.002902497,
  0, -0.01376272, -0.00969515, -0.004411527, -0.0007787212, 0.0007787212, 
    0.004411527, 0.00969515, 0.01376272, 0,
  0, 0.001673691, -0.008278607, -0.006019558, -0.00200568, 0.00200568, 
    0.006019558, 0.008278607, -0.001673691, 0,
  0, 0, -0.000388854, -0.002758372, -0.0005684611, 0.0005684611, 0.002758372, 
    0.000388854, 0, 0,
  0, 0, 0, 0, 0.0001421608, -0.0001421608, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0001378467, -0.0001378467, 0, 0, 0, 0,
  0, 0, -0.0002449594, -0.002685626, -0.0005441869, 0.0005441869, 
    0.002685626, 0.0002449594, 0, 0,
  0, 0.00179794, -0.008016966, -0.005816287, -0.001922676, 0.001922676, 
    0.005816287, 0.008016966, -0.00179794, 0,
  0, -0.01334754, -0.009357425, -0.004169604, -0.0007107307, 0.0007107307, 
    0.004169604, 0.009357425, 0.01334754, 0,
  0.002811883, -0.01051145, -0.0102144, -0.002035744, -0.0001187086, 
    0.0001187086, 0.002035744, 0.0102144, 0.01051145, -0.002811883,
  0.002811883, -0.01051145, -0.0102144, -0.002035744, -0.0001187086, 
    0.0001187086, 0.002035744, 0.0102144, 0.01051145, -0.002811883,
  0, -0.01334754, -0.009357425, -0.004169604, -0.0007107307, 0.0007107307, 
    0.004169604, 0.009357425, 0.01334754, 0,
  0, 0.00179794, -0.008016966, -0.005816287, -0.001922676, 0.001922676, 
    0.005816287, 0.008016966, -0.00179794, 0,
  0, 0, -0.0002449594, -0.002685626, -0.0005441869, 0.0005441869, 
    0.002685626, 0.0002449594, 0, 0,
  0, 0, 0, 0, 0.0001378467, -0.0001378467, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0001258095, -0.0001258095, 0, 0, 0, 0,
  0, 0, -0.0001249876, -0.002491703, -0.0004913866, 0.0004913866, 
    0.002491703, 0.0001249876, 0, 0,
  0, 0.001794341, -0.007418247, -0.005371028, -0.001767041, 0.001767041, 
    0.005371028, 0.007418247, -0.001794341, 0,
  0, -0.01234152, -0.008632522, -0.003793863, -0.0006244552, 0.0006244552, 
    0.003793863, 0.008632522, 0.01234152, 0,
  0.002593941, -0.009686967, -0.009397025, -0.001792832, -0.0001002306, 
    0.0001002306, 0.001792832, 0.009397025, 0.009686967, -0.002593941,
  0.002593941, -0.009686967, -0.009397025, -0.001792832, -0.0001002306, 
    0.0001002306, 0.001792832, 0.009397025, 0.009686967, -0.002593941,
  0, -0.01234152, -0.008632522, -0.003793863, -0.0006244552, 0.0006244552, 
    0.003793863, 0.008632522, 0.01234152, 0,
  0, 0.001794341, -0.007418247, -0.005371028, -0.001767041, 0.001767041, 
    0.005371028, 0.007418247, -0.001794341, 0,
  0, 0, -0.0001249876, -0.002491703, -0.0004913866, 0.0004913866, 
    0.002491703, 0.0001249876, 0, 0,
  0, 0, 0, 0, 0.0001258095, -0.0001258095, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0001080338, -0.0001080338, 0, 0, 0, 0,
  0, 0, -4.305307e-05, -0.002182445, -0.0004181444, 0.0004181444, 
    0.002182445, 4.305307e-05, 0, 0,
  0, 0.00165294, -0.006489325, -0.00469028, -0.001540245, 0.001540245, 
    0.00469028, 0.006489325, -0.00165294, 0,
  0, -0.01078118, -0.007531179, -0.003285282, -0.000527743, 0.000527743, 
    0.003285282, 0.007531179, 0.01078118, 0,
  0.002259423, -0.008433656, -0.008196944, -0.00151723, -8.128507e-05, 
    8.128507e-05, 0.00151723, 0.008196944, 0.008433656, -0.002259423,
  0.002259423, -0.008433656, -0.008196944, -0.00151723, -8.128507e-05, 
    8.128507e-05, 0.00151723, 0.008196944, 0.008433656, -0.002259423,
  0, -0.01078118, -0.007531179, -0.003285282, -0.000527743, 0.000527743, 
    0.003285282, 0.007531179, 0.01078118, 0,
  0, 0.00165294, -0.006489325, -0.00469028, -0.001540245, 0.001540245, 
    0.00469028, 0.006489325, -0.00165294, 0,
  0, 0, -4.305307e-05, -0.002182445, -0.0004181444, 0.0004181444, 
    0.002182445, 4.305307e-05, 0, 0,
  0, 0, 0, 0, 0.0001080338, -0.0001080338, 0, 0, 0, 0,
  0, 0, 0, 0, 8.704685e-05, -8.704685e-05, 0, 0, 0, 0,
  0, 0, 6.148277e-06, -0.001792324, -0.0003342622, 0.0003342622, 0.001792324, 
    -6.148277e-06, 0, 0,
  0, 0.00140789, -0.005325592, -0.003842935, -0.001261296, 0.001261296, 
    0.003842935, 0.005325592, -0.00140789, 0,
  0, -0.008835113, -0.006165193, -0.00267771, -0.0004233849, 0.0004233849, 
    0.00267771, 0.006165193, 0.008835113, 0,
  0.00184585, -0.006888379, -0.006716882, -0.001217658, -6.336612e-05, 
    6.336612e-05, 0.001217658, 0.006716882, 0.006888379, -0.00184585,
  0.00184585, -0.006888379, -0.006716882, -0.001217658, -6.336612e-05, 
    6.336612e-05, 0.001217658, 0.006716882, 0.006888379, -0.00184585,
  0, -0.008835113, -0.006165193, -0.00267771, -0.0004233849, 0.0004233849, 
    0.00267771, 0.006165193, 0.008835113, 0,
  0, 0.00140789, -0.005325592, -0.003842935, -0.001261296, 0.001261296, 
    0.003842935, 0.005325592, -0.00140789, 0,
  0, 0, 6.148277e-06, -0.001792324, -0.0003342622, 0.0003342622, 0.001792324, 
    -6.148277e-06, 0, 0,
  0, 0, 0, 0, 8.704685e-05, -8.704685e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 6.474754e-05, -6.474754e-05, 0, 0, 0, 0,
  0, 0, 2.915298e-05, -0.001356237, -0.0002468703, 0.0002468703, 0.001356237, 
    -2.915298e-05, 0, 0,
  0, 0.001094844, -0.004027885, -0.002901813, -0.0009523921, 0.0009523921, 
    0.002901813, 0.004027885, -0.001094844, 0,
  0, -0.006673533, -0.004651777, -0.002014543, -0.0003151065, 0.0003151065, 
    0.002014543, 0.004651777, 0.006673533, 0,
  0.001389731, -0.005185776, -0.005074942, -0.0009061344, -4.640701e-05, 
    4.640701e-05, 0.0009061344, 0.005074942, 0.005185776, -0.001389731,
  0.001389731, -0.005185776, -0.005074942, -0.0009061344, -4.640701e-05, 
    4.640701e-05, 0.0009061344, 0.005074942, 0.005185776, -0.001389731,
  0, -0.006673533, -0.004651777, -0.002014543, -0.0003151065, 0.0003151065, 
    0.002014543, 0.004651777, 0.006673533, 0,
  0, 0.001094844, -0.004027885, -0.002901813, -0.0009523921, 0.0009523921, 
    0.002901813, 0.004027885, -0.001094844, 0,
  0, 0, 2.915298e-05, -0.001356237, -0.0002468703, 0.0002468703, 0.001356237, 
    -2.915298e-05, 0, 0,
  0, 0, 0, 0, 6.474754e-05, -6.474754e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 4.238164e-05, -4.238164e-05, 0, 0, 0, 0,
  0, 0, 3.225733e-05, -0.0009015123, -0.0001605106, 0.0001605106, 
    0.0009015123, -3.225733e-05, 0, 0,
  0, 0.0007430961, -0.002676153, -0.001924598, -0.0006317715, 0.0006317715, 
    0.001924598, 0.002676153, -0.0007430961, 0,
  0, -0.004429145, -0.00308317, -0.001332187, -0.0002067488, 0.0002067488, 
    0.001332187, 0.00308317, 0.004429145, 0,
  0.0009189562, -0.003429061, -0.003368417, -0.0005942997, -3.021932e-05, 
    3.021932e-05, 0.0005942997, 0.003368417, 0.003429061, -0.0009189562,
  0.0009189562, -0.003429061, -0.003368417, -0.0005942997, -3.021932e-05, 
    3.021932e-05, 0.0005942997, 0.003368417, 0.003429061, -0.0009189562,
  0, -0.004429145, -0.00308317, -0.001332187, -0.0002067488, 0.0002067488, 
    0.001332187, 0.00308317, 0.004429145, 0,
  0, 0.0007430961, -0.002676153, -0.001924598, -0.0006317715, 0.0006317715, 
    0.001924598, 0.002676153, -0.0007430961, 0,
  0, 0, 3.225733e-05, -0.0009015123, -0.0001605106, 0.0001605106, 
    0.0009015123, -3.225733e-05, 0, 0,
  0, 0, 0, 0, 4.238164e-05, -4.238164e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 2.069441e-05, -2.069441e-05, 0, 0, 0, 0,
  0, 0, 2.117404e-05, -0.0004464598, -7.782724e-05, 7.782724e-05, 
    0.0004464598, -2.117404e-05, 0, 0,
  0, 0.0003742031, -0.001324471, -0.0009508296, -0.000312237, 0.000312237, 
    0.0009508296, 0.001324471, -0.0003742031, 0,
  0, -0.00219062, -0.001522253, -0.0006564604, -0.0001012366, 0.0001012366, 
    0.0006564604, 0.001522253, 0.00219062, 0,
  0.0004523387, -0.001687976, -0.001665744, -0.0002908438, -1.477318e-05, 
    1.477318e-05, 0.0002908438, 0.001665744, 0.001687976, -0.0004523387,
  0.0004523387, -0.001687976, -0.001665744, -0.0002908438, -1.477318e-05, 
    1.477318e-05, 0.0002908438, 0.001665744, 0.001687976, -0.0004523387,
  0, -0.00219062, -0.001522253, -0.0006564604, -0.0001012366, 0.0001012366, 
    0.0006564604, 0.001522253, 0.00219062, 0,
  0, 0.0003742031, -0.001324471, -0.0009508296, -0.000312237, 0.000312237, 
    0.0009508296, 0.001324471, -0.0003742031, 0,
  0, 0, 2.117404e-05, -0.0004464598, -7.782724e-05, 7.782724e-05, 
    0.0004464598, -2.117404e-05, 0, 0,
  0, 0, 0, 0, 2.069441e-05, -2.069441e-05, 0, 0, 0, 0,
  0, 0, 0, 0, -3.793572e-10, 3.793572e-10, 0, 0, 0, 0,
  0, 0, -1.268874e-08, -6.309733e-09, -2.031081e-09, 2.031081e-09, 
    6.309733e-09, 1.268874e-08, 0, 0,
  0, -1.176477e-08, -2.342423e-08, -1.542942e-08, -4.979319e-09, 
    4.979319e-09, 1.542942e-08, 2.342423e-08, 1.176477e-08, 0,
  0, -3.397442e-08, -2.524942e-08, -1.542458e-08, -5.082796e-09, 
    5.082796e-09, 1.542458e-08, 2.524942e-08, 3.397442e-08, 0,
  8.218023e-09, -3.649568e-08, -2.59674e-08, -1.529537e-08, -5.735643e-09, 
    5.735643e-09, 1.529537e-08, 2.59674e-08, 3.649568e-08, -8.218023e-09,
  8.218023e-09, -3.649568e-08, -2.59674e-08, -1.529537e-08, -5.735643e-09, 
    5.735643e-09, 1.529537e-08, 2.59674e-08, 3.649568e-08, -8.218023e-09,
  0, -3.397442e-08, -2.524942e-08, -1.542458e-08, -5.082796e-09, 
    5.082796e-09, 1.542458e-08, 2.524942e-08, 3.397442e-08, 0,
  0, -1.176477e-08, -2.342423e-08, -1.542942e-08, -4.979319e-09, 
    4.979319e-09, 1.542942e-08, 2.342423e-08, 1.176477e-08, 0,
  0, 0, -1.268874e-08, -6.309733e-09, -2.031081e-09, 2.031081e-09, 
    6.309733e-09, 1.268874e-08, 0, 0,
  0, 0, 0, 0, -3.793572e-10, 3.793572e-10, 0, 0, 0, 0,
  0, 0, 0, 2.937466e-05, 2.721521e-05, -2.721521e-05, -2.937466e-05, 0, 0, 0,
  0, 0, -0.0002436649, -0.0001216534, -0.0001020982, 0.0001020982, 
    0.0001216534, 0.0002436649, 0, 0,
  0, -0.0006781258, -0.00828121, -0.005612711, -0.001733972, 0.001733972, 
    0.005612711, 0.00828121, 0.0006781258, 0,
  0.0005927979, -0.002210401, -0.009385014, -0.004610501, -0.0008418286, 
    0.0008418286, 0.004610501, 0.009385014, 0.002210401, -0.0005927979,
  0.0009220587, -0.003447537, -0.009744491, -0.002375761, -0.000137582, 
    0.000137582, 0.002375761, 0.009744491, 0.003447537, -0.0009220587,
  0.0009220587, -0.003447537, -0.009744491, -0.002375761, -0.000137582, 
    0.000137582, 0.002375761, 0.009744491, 0.003447537, -0.0009220587,
  0.0005927979, -0.002210401, -0.009385014, -0.004610501, -0.0008418286, 
    0.0008418286, 0.004610501, 0.009385014, 0.002210401, -0.0005927979,
  0, -0.0006781258, -0.00828121, -0.005612711, -0.001733972, 0.001733972, 
    0.005612711, 0.00828121, 0.0006781258, 0,
  0, 0, -0.0002436649, -0.0001216534, -0.0001020982, 0.0001020982, 
    0.0001216534, 0.0002436649, 0, 0,
  0, 0, 0, 2.937466e-05, 2.721521e-05, -2.721521e-05, -2.937466e-05, 0, 0, 0,
  0, 0, 0, 2.753662e-05, 2.698793e-05, -2.698793e-05, -2.753662e-05, 0, 0, 0,
  0, 0, -0.0001997186, -0.0001145652, -0.000101137, 0.000101137, 
    0.0001145652, 0.0001997186, 0, 0,
  0, -0.0006111048, -0.008210798, -0.005550113, -0.001709998, 0.001709998, 
    0.005550113, 0.008210798, 0.0006111048, 0,
  0.0005801168, -0.002162982, -0.009281811, -0.00453299, -0.0008118864, 
    0.0008118864, 0.00453299, 0.009281811, 0.002162982, -0.0005801168,
  0.0009105077, -0.00340015, -0.009612685, -0.002300074, -0.0001294365, 
    0.0001294365, 0.002300074, 0.009612685, 0.00340015, -0.0009105077,
  0.0009105077, -0.00340015, -0.009612685, -0.002300074, -0.0001294365, 
    0.0001294365, 0.002300074, 0.009612685, 0.00340015, -0.0009105077,
  0.0005801168, -0.002162982, -0.009281811, -0.00453299, -0.0008118864, 
    0.0008118864, 0.00453299, 0.009281811, 0.002162982, -0.0005801168,
  0, -0.0006111048, -0.008210798, -0.005550113, -0.001709998, 0.001709998, 
    0.005550113, 0.008210798, 0.0006111048, 0,
  0, 0, -0.0001997186, -0.0001145652, -0.000101137, 0.000101137, 
    0.0001145652, 0.0001997186, 0, 0,
  0, 0, 0, 2.753662e-05, 2.698793e-05, -2.698793e-05, -2.753662e-05, 0, 0, 0,
  0, 0, 0, 2.459871e-05, 2.619718e-05, -2.619718e-05, -2.459871e-05, 0, 0, 0,
  0, 0, -0.0001212417, -0.0001018609, -9.80252e-05, 9.80252e-05, 
    0.0001018609, 0.0001212417, 0, 0,
  0, -0.0004923516, -0.007942389, -0.005351122, -0.001640004, 0.001640004, 
    0.005351122, 0.007942389, 0.0004923516, 0,
  0.0005478773, -0.002043155, -0.008962078, -0.004296739, -0.0007429817, 
    0.0007429817, 0.004296739, 0.008962078, 0.002043155, -0.0005478773,
  0.0008747906, -0.003264622, -0.009233337, -0.00210894, -0.0001134368, 
    0.0001134368, 0.00210894, 0.009233337, 0.003264622, -0.0008747906,
  0.0008747906, -0.003264622, -0.009233337, -0.00210894, -0.0001134368, 
    0.0001134368, 0.00210894, 0.009233337, 0.003264622, -0.0008747906,
  0.0005478773, -0.002043155, -0.008962078, -0.004296739, -0.0007429817, 
    0.0007429817, 0.004296739, 0.008962078, 0.002043155, -0.0005478773,
  0, -0.0004923516, -0.007942389, -0.005351122, -0.001640004, 0.001640004, 
    0.005351122, 0.007942389, 0.0004923516, 0,
  0, 0, -0.0001212417, -0.0001018609, -9.80252e-05, 9.80252e-05, 
    0.0001018609, 0.0001212417, 0, 0,
  0, 0, 0, 2.459871e-05, 2.619718e-05, -2.619718e-05, -2.459871e-05, 0, 0, 0,
  0, 0, 0, 2.114013e-05, 2.395063e-05, -2.395063e-05, -2.114013e-05, 0, 0, 0,
  0, 0, -5.588763e-05, -8.658683e-05, -8.959212e-05, 8.959212e-05, 
    8.658683e-05, 5.588763e-05, 0, 0,
  0, -0.0003777269, -0.007337223, -0.004942738, -0.001511542, 0.001511542, 
    0.004942738, 0.007337223, 0.0003777269, 0,
  0.0004952688, -0.001847067, -0.008294187, -0.003911743, -0.0006553119, 
    0.0006553119, 0.003911743, 0.008294187, 0.001847067, -0.0004952688,
  0.0008008862, -0.002988057, -0.008522817, -0.001860625, -9.445607e-05, 
    9.445607e-05, 0.001860625, 0.008522817, 0.002988057, -0.0008008862,
  0.0008008862, -0.002988057, -0.008522817, -0.001860625, -9.445607e-05, 
    9.445607e-05, 0.001860625, 0.008522817, 0.002988057, -0.0008008862,
  0.0004952688, -0.001847067, -0.008294187, -0.003911743, -0.0006553119, 
    0.0006553119, 0.003911743, 0.008294187, 0.001847067, -0.0004952688,
  0, -0.0003777269, -0.007337223, -0.004942738, -0.001511542, 0.001511542, 
    0.004942738, 0.007337223, 0.0003777269, 0,
  0, 0, -5.588763e-05, -8.658683e-05, -8.959212e-05, 8.959212e-05, 
    8.658683e-05, 5.588763e-05, 0, 0,
  0, 0, 0, 2.114013e-05, 2.395063e-05, -2.395063e-05, -2.114013e-05, 0, 0, 0,
  0, 0, 0, 1.734022e-05, 2.057202e-05, -2.057202e-05, -1.734022e-05, 0, 0, 0,
  0, 0, -1.112143e-05, -7.011503e-05, -7.694183e-05, 7.694183e-05, 
    7.011503e-05, 1.112143e-05, 0, 0,
  0, -0.0002782268, -0.006408261, -0.004321288, -0.001321844, 0.001321844, 
    0.004321288, 0.006408261, 0.0002782268, 0,
  0.0004246696, -0.001583891, -0.007265355, -0.003385333, -0.0005555307, 
    0.0005555307, 0.003385333, 0.007265355, 0.001583891, -0.0004246696,
  0.0006926283, -0.002583976, -0.007463949, -0.001574976, -7.596873e-05, 
    7.596873e-05, 0.001574976, 0.007463949, 0.002583976, -0.0006926283,
  0.0006926283, -0.002583976, -0.007463949, -0.001574976, -7.596873e-05, 
    7.596873e-05, 0.001574976, 0.007463949, 0.002583976, -0.0006926283,
  0.0004246696, -0.001583891, -0.007265355, -0.003385333, -0.0005555307, 
    0.0005555307, 0.003385333, 0.007265355, 0.001583891, -0.0004246696,
  0, -0.0002782268, -0.006408261, -0.004321288, -0.001321844, 0.001321844, 
    0.004321288, 0.006408261, 0.0002782268, 0,
  0, 0, -1.112143e-05, -7.011503e-05, -7.694183e-05, 7.694183e-05, 
    7.011503e-05, 1.112143e-05, 0, 0,
  0, 0, 0, 1.734022e-05, 2.057202e-05, -2.057202e-05, -1.734022e-05, 0, 0, 0,
  0, 0, 0, 1.346958e-05, 1.65724e-05, -1.65724e-05, -1.346958e-05, 0, 0, 0,
  0, 0, 1.515912e-05, -5.373624e-05, -6.196715e-05, 6.196715e-05, 
    5.373624e-05, -1.515912e-05, 0, 0,
  0, -0.0001949756, -0.005252321, -0.003545666, -0.001085737, 0.001085737, 
    0.003545666, 0.005252321, 0.0001949756, 0,
  0.0003426427, -0.001278079, -0.00597164, -0.00275675, -0.0004466841, 
    0.0004466841, 0.00275675, 0.00597164, 0.001278079, -0.0003426427,
  0.0005622989, -0.002097788, -0.006139196, -0.001263427, -5.899592e-05, 
    5.899592e-05, 0.001263427, 0.006139196, 0.002097788, -0.0005622989,
  0.0005622989, -0.002097788, -0.006139196, -0.001263427, -5.899592e-05, 
    5.899592e-05, 0.001263427, 0.006139196, 0.002097788, -0.0005622989,
  0.0003426427, -0.001278079, -0.00597164, -0.00275675, -0.0004466841, 
    0.0004466841, 0.00275675, 0.00597164, 0.001278079, -0.0003426427,
  0, -0.0001949756, -0.005252321, -0.003545666, -0.001085737, 0.001085737, 
    0.003545666, 0.005252321, 0.0001949756, 0,
  0, 0, 1.515912e-05, -5.373624e-05, -6.196715e-05, 6.196715e-05, 
    5.373624e-05, -1.515912e-05, 0, 0,
  0, 0, 0, 1.346958e-05, 1.65724e-05, -1.65724e-05, -1.346958e-05, 0, 0, 0,
  0, 0, 0, 9.73296e-06, 1.231937e-05, -1.231937e-05, -9.73296e-06, 0, 0, 0,
  0, 0, 2.597713e-05, -3.829425e-05, -4.604799e-05, 4.604799e-05, 
    3.829425e-05, -2.597713e-05, 0, 0,
  0, -0.0001277715, -0.003969084, -0.002681595, -0.0008220871, 0.0008220871, 
    0.002681595, 0.003969084, 0.0001277715, 0,
  0.0002554594, -0.0009529833, -0.004523174, -0.002072225, -0.0003330655, 
    0.0003330655, 0.002072225, 0.004523174, 0.0009529833, -0.0002554594,
  0.0004210924, -0.001571069, -0.004654329, -0.000939663, -4.315929e-05, 
    4.315929e-05, 0.000939663, 0.004654329, 0.001571069, -0.0004210924,
  0.0004210924, -0.001571069, -0.004654329, -0.000939663, -4.315929e-05, 
    4.315929e-05, 0.000939663, 0.004654329, 0.001571069, -0.0004210924,
  0.0002554594, -0.0009529833, -0.004523174, -0.002072225, -0.0003330655, 
    0.0003330655, 0.002072225, 0.004523174, 0.0009529833, -0.0002554594,
  0, -0.0001277715, -0.003969084, -0.002681595, -0.0008220871, 0.0008220871, 
    0.002681595, 0.003969084, 0.0001277715, 0,
  0, 0, 2.597713e-05, -3.829425e-05, -4.604799e-05, 4.604799e-05, 
    3.829425e-05, -2.597713e-05, 0, 0,
  0, 0, 0, 9.73296e-06, 1.231937e-05, -1.231937e-05, -9.73296e-06, 0, 0, 0,
  0, 0, 0, 6.229418e-06, 8.053987e-06, -8.053987e-06, -6.229418e-06, 0, 0, 0,
  0, 0, 2.485497e-05, -2.415505e-05, -3.009092e-05, 3.009092e-05, 
    2.415505e-05, -2.485497e-05, 0, 0,
  0, -7.482824e-05, -0.002636307, -0.001781949, -0.0005467999, 0.0005467999, 
    0.001781949, 0.002636307, 7.482824e-05, 0,
  0.0001676652, -0.000625542, -0.003009646, -0.001369582, -0.0002189408, 
    0.0002189408, 0.001369582, 0.003009646, 0.000625542, -0.0001676652,
  0.0002771921, -0.001034266, -0.003099435, -0.0006161059, -2.812003e-05, 
    2.812003e-05, 0.0006161059, 0.003099435, 0.001034266, -0.0002771921,
  0.0002771921, -0.001034266, -0.003099435, -0.0006161059, -2.812003e-05, 
    2.812003e-05, 0.0006161059, 0.003099435, 0.001034266, -0.0002771921,
  0.0001676652, -0.000625542, -0.003009646, -0.001369582, -0.0002189408, 
    0.0002189408, 0.001369582, 0.003009646, 0.000625542, -0.0001676652,
  0, -7.482824e-05, -0.002636307, -0.001781949, -0.0005467999, 0.0005467999, 
    0.001781949, 0.002636307, 7.482824e-05, 0,
  0, 0, 2.485497e-05, -2.415505e-05, -3.009092e-05, 3.009092e-05, 
    2.415505e-05, -2.485497e-05, 0, 0,
  0, 0, 0, 6.229418e-06, 8.053987e-06, -8.053987e-06, -6.229418e-06, 0, 0, 0,
  0, 0, 0, 2.978258e-06, 3.9232e-06, -3.9232e-06, -2.978258e-06, 0, 0, 0,
  0, 0, 1.538461e-05, -1.13621e-05, -1.464857e-05, 1.464857e-05, 1.13621e-05, 
    -1.538461e-05, 0, 0,
  0, -3.311473e-05, -0.00130512, -0.000882685, -0.0002710968, 0.0002710968, 
    0.000882685, 0.00130512, 3.311473e-05, 0,
  8.20508e-05, -0.0003061637, -0.00149255, -0.0006751646, -0.000107478, 
    0.000107478, 0.0006751646, 0.00149255, 0.0003061637, -8.20508e-05,
  0.0001358988, -0.0005071203, -0.00153842, -0.0003017059, -1.377299e-05, 
    1.377299e-05, 0.0003017059, 0.00153842, 0.0005071203, -0.0001358988,
  0.0001358988, -0.0005071203, -0.00153842, -0.0003017059, -1.377299e-05, 
    1.377299e-05, 0.0003017059, 0.00153842, 0.0005071203, -0.0001358988,
  8.20508e-05, -0.0003061637, -0.00149255, -0.0006751646, -0.000107478, 
    0.000107478, 0.0006751646, 0.00149255, 0.0003061637, -8.20508e-05,
  0, -3.311473e-05, -0.00130512, -0.000882685, -0.0002710968, 0.0002710968, 
    0.000882685, 0.00130512, 3.311473e-05, 0,
  0, 0, 1.538461e-05, -1.13621e-05, -1.464857e-05, 1.464857e-05, 1.13621e-05, 
    -1.538461e-05, 0, 0,
  0, 0, 0, 2.978258e-06, 3.9232e-06, -3.9232e-06, -2.978258e-06, 0, 0, 0,
  0, 0, 0, 5.853413e-10, 3.118638e-10, -3.118638e-10, -5.853413e-10, 0, 0, 0,
  0, 0, -1.151457e-08, -4.234781e-09, -1.096469e-09, 1.096469e-09, 
    4.234781e-09, 1.151457e-08, 0, 0,
  0, -1.320141e-08, -2.347333e-08, -1.558718e-08, -4.875147e-09, 
    4.875147e-09, 1.558718e-08, 2.347333e-08, 1.320141e-08, 0,
  5.808732e-09, -2.375368e-08, -2.46941e-08, -1.544228e-08, -5.093391e-09, 
    5.093391e-09, 1.544228e-08, 2.46941e-08, 2.375368e-08, -5.808732e-09,
  7.001435e-09, -2.863566e-08, -2.551781e-08, -1.530671e-08, -5.799936e-09, 
    5.799936e-09, 1.530671e-08, 2.551781e-08, 2.863566e-08, -7.001435e-09,
  7.001435e-09, -2.863566e-08, -2.551781e-08, -1.530671e-08, -5.799936e-09, 
    5.799936e-09, 1.530671e-08, 2.551781e-08, 2.863566e-08, -7.001435e-09,
  5.808732e-09, -2.375368e-08, -2.46941e-08, -1.544228e-08, -5.093391e-09, 
    5.093391e-09, 1.544228e-08, 2.46941e-08, 2.375368e-08, -5.808732e-09,
  0, -1.320141e-08, -2.347333e-08, -1.558718e-08, -4.875147e-09, 
    4.875147e-09, 1.558718e-08, 2.347333e-08, 1.320141e-08, 0,
  0, 0, -1.151457e-08, -4.234781e-09, -1.096469e-09, 1.096469e-09, 
    4.234781e-09, 1.151457e-08, 0, 0,
  0, 0, 0, 5.853413e-10, 3.118638e-10, -3.118638e-10, -5.853413e-10, 0, 0, 0,
  0, 0, 0, 3.046667e-05, 2.745757e-05, -2.745757e-05, -3.046667e-05, 0, 0, 0,
  0, 0, -0.0002546235, -0.0001257831, -0.00010299, 0.00010299, 0.0001257831, 
    0.0002546235, 0, 0,
  0, -0.0006940318, -0.00828829, -0.005597732, -0.001725802, 0.001725802, 
    0.005597732, 0.00828829, 0.0006940318, 0,
  0.0005976551, -0.002228644, -0.009351598, -0.004594702, -0.0008440774, 
    0.0008440774, 0.004594702, 0.009351598, 0.002228644, -0.0005976551,
  0.0009266008, -0.00346467, -0.009684209, -0.002380941, -0.0001401419, 
    0.0001401419, 0.002380941, 0.009684209, 0.00346467, -0.0009266008,
  0.0009266008, -0.00346467, -0.009684209, -0.002380941, -0.0001401419, 
    0.0001401419, 0.002380941, 0.009684209, 0.00346467, -0.0009266008,
  0.0005976551, -0.002228644, -0.009351598, -0.004594702, -0.0008440774, 
    0.0008440774, 0.004594702, 0.009351598, 0.002228644, -0.0005976551,
  0, -0.0006940318, -0.00828829, -0.005597732, -0.001725802, 0.001725802, 
    0.005597732, 0.00828829, 0.0006940318, 0,
  0, 0, -0.0002546235, -0.0001257831, -0.00010299, 0.00010299, 0.0001257831, 
    0.0002546235, 0, 0,
  0, 0, 0, 3.046667e-05, 2.745757e-05, -2.745757e-05, -3.046667e-05, 0, 0, 0,
  0, 0, 0, 2.863302e-05, 2.72283e-05, -2.72283e-05, -2.863302e-05, 0, 0, 0,
  0, 0, -0.0002107615, -0.0001186984, -0.0001020216, 0.0001020216, 
    0.0001186984, 0.0002107615, 0, 0,
  0, -0.0006271242, -0.008217847, -0.005535415, -0.001702062, 0.001702062, 
    0.005535415, 0.008217847, 0.0006271242, 0,
  0.000584978, -0.002181178, -0.00924895, -0.004517405, -0.0008142332, 
    0.0008142332, 0.004517405, 0.00924895, 0.002181178, -0.000584978,
  0.0009150683, -0.003417269, -0.009553849, -0.002305315, -0.0001318761, 
    0.0001318761, 0.002305315, 0.009553849, 0.003417269, -0.0009150683,
  0.0009150683, -0.003417269, -0.009553849, -0.002305315, -0.0001318761, 
    0.0001318761, 0.002305315, 0.009553849, 0.003417269, -0.0009150683,
  0.000584978, -0.002181178, -0.00924895, -0.004517405, -0.0008142332, 
    0.0008142332, 0.004517405, 0.00924895, 0.002181178, -0.000584978,
  0, -0.0006271242, -0.008217847, -0.005535415, -0.001702062, 0.001702062, 
    0.005535415, 0.008217847, 0.0006271242, 0,
  0, 0, -0.0002107615, -0.0001186984, -0.0001020216, 0.0001020216, 
    0.0001186984, 0.0002107615, 0, 0,
  0, 0, 0, 2.863302e-05, 2.72283e-05, -2.72283e-05, -2.863302e-05, 0, 0, 0,
  0, 0, 0, 2.568198e-05, 2.642871e-05, -2.642871e-05, -2.568198e-05, 0, 0, 0,
  0, 0, -0.0001321262, -0.0001059302, -9.887929e-05, 9.887929e-05, 
    0.0001059302, 0.0001321262, 0, 0,
  0, -0.0005080745, -0.007949643, -0.005337188, -0.001632569, 0.001632569, 
    0.005337188, 0.007949643, 0.0005080745, 0,
  0.0005526862, -0.002061121, -0.008930719, -0.004282035, -0.000745484, 
    0.000745484, 0.004282035, 0.008930719, 0.002061121, -0.0005526862,
  0.0008792863, -0.00328145, -0.009177702, -0.002114474, -0.000115579, 
    0.000115579, 0.002114474, 0.009177702, 0.00328145, -0.0008792863,
  0.0008792863, -0.00328145, -0.009177702, -0.002114474, -0.000115579, 
    0.000115579, 0.002114474, 0.009177702, 0.00328145, -0.0008792863,
  0.0005526862, -0.002061121, -0.008930719, -0.004282035, -0.000745484, 
    0.000745484, 0.004282035, 0.008930719, 0.002061121, -0.0005526862,
  0, -0.0005080745, -0.007949643, -0.005337188, -0.001632569, 0.001632569, 
    0.005337188, 0.007949643, 0.0005080745, 0,
  0, 0, -0.0001321262, -0.0001059302, -9.887929e-05, 9.887929e-05, 
    0.0001059302, 0.0001321262, 0, 0,
  0, 0, 0, 2.568198e-05, 2.642871e-05, -2.642871e-05, -2.568198e-05, 0, 0, 0,
  0, 0, 0, 2.215118e-05, 2.416347e-05, -2.416347e-05, -2.215118e-05, 0, 0, 0,
  0, 0, -6.606273e-05, -9.037773e-05, -9.037944e-05, 9.037944e-05, 
    9.037773e-05, 6.606273e-05, 0, 0,
  0, -0.0003924186, -0.007344917, -0.004930267, -0.001504841, 0.001504841, 
    0.004930267, 0.007344917, 0.0003924186, 0,
  0.0004998034, -0.001863993, -0.008265833, -0.00389852, -0.0006578621, 
    0.0006578621, 0.00389852, 0.008265833, 0.001863993, -0.0004998034,
  0.0008051077, -0.003003838, -0.0084723, -0.00186627, -9.625436e-05, 
    9.625436e-05, 0.00186627, 0.0084723, 0.003003838, -0.0008051077,
  0.0008051077, -0.003003838, -0.0084723, -0.00186627, -9.625436e-05, 
    9.625436e-05, 0.00186627, 0.0084723, 0.003003838, -0.0008051077,
  0.0004998034, -0.001863993, -0.008265833, -0.00389852, -0.0006578621, 
    0.0006578621, 0.00389852, 0.008265833, 0.001863993, -0.0004998034,
  0, -0.0003924186, -0.007344917, -0.004930267, -0.001504841, 0.001504841, 
    0.004930267, 0.007344917, 0.0003924186, 0,
  0, 0, -6.606273e-05, -9.037773e-05, -9.037944e-05, 9.037944e-05, 
    9.037773e-05, 6.606273e-05, 0, 0,
  0, 0, 0, 2.215118e-05, 2.416347e-05, -2.416347e-05, -2.215118e-05, 0, 0, 0,
  0, 0, 0, 1.822705e-05, 2.07577e-05, -2.07577e-05, -1.822705e-05, 0, 0, 0,
  0, 0, -2.007348e-05, -7.34364e-05, -7.763013e-05, 7.763013e-05, 
    7.34364e-05, 2.007348e-05, 0, 0,
  0, -0.0002912104, -0.006416466, -0.00431102, -0.001316148, 0.001316148, 
    0.00431102, 0.006416466, 0.0002912104, 0,
  0.0004287128, -0.001598977, -0.007241611, -0.00337412, -0.0005579437, 
    0.0005579437, 0.00337412, 0.007241611, 0.001598977, -0.0004287128,
  0.0006963831, -0.002598002, -0.007420705, -0.001580322, -7.744075e-05, 
    7.744075e-05, 0.001580322, 0.007420705, 0.002598002, -0.0006963831,
  0.0006963831, -0.002598002, -0.007420705, -0.001580322, -7.744075e-05, 
    7.744075e-05, 0.001580322, 0.007420705, 0.002598002, -0.0006963831,
  0.0004287128, -0.001598977, -0.007241611, -0.00337412, -0.0005579437, 
    0.0005579437, 0.00337412, 0.007241611, 0.001598977, -0.0004287128,
  0, -0.0002912104, -0.006416466, -0.00431102, -0.001316148, 0.001316148, 
    0.00431102, 0.006416466, 0.0002912104, 0,
  0, 0, -2.007348e-05, -7.34364e-05, -7.763013e-05, 7.763013e-05, 
    7.34364e-05, 2.007348e-05, 0, 0,
  0, 0, 0, 1.822705e-05, 2.07577e-05, -2.07577e-05, -1.822705e-05, 0, 0, 0,
  0, 0, 0, 1.419874e-05, 1.672446e-05, -1.672446e-05, -1.419874e-05, 0, 0, 0,
  0, 0, 7.749403e-06, -5.646477e-05, -6.253186e-05, 6.253186e-05, 
    5.646477e-05, -7.749403e-06, 0, 0,
  0, -0.0002058307, -0.005260962, -0.003538133, -0.001081273, 0.001081273, 
    0.003538133, 0.005260962, 0.0002058307, 0,
  0.0003460448, -0.001290771, -0.005953672, -0.002747942, -0.000448809, 
    0.000448809, 0.002747942, 0.005953672, 0.001290771, -0.0003460448,
  0.0005654459, -0.002109539, -0.006104944, -0.001268135, -6.016145e-05, 
    6.016145e-05, 0.001268135, 0.006104944, 0.002109539, -0.0005654459,
  0.0005654459, -0.002109539, -0.006104944, -0.001268135, -6.016145e-05, 
    6.016145e-05, 0.001268135, 0.006104944, 0.002109539, -0.0005654459,
  0.0003460448, -0.001290771, -0.005953672, -0.002747942, -0.000448809, 
    0.000448809, 0.002747942, 0.005953672, 0.001290771, -0.0003460448,
  0, -0.0002058307, -0.005260962, -0.003538133, -0.001081273, 0.001081273, 
    0.003538133, 0.005260962, 0.0002058307, 0,
  0, 0, 7.749403e-06, -5.646477e-05, -6.253186e-05, 6.253186e-05, 
    5.646477e-05, -7.749403e-06, 0, 0,
  0, 0, 0, 1.419874e-05, 1.672446e-05, -1.672446e-05, -1.419874e-05, 0, 0, 0,
  0, 0, 0, 1.02857e-05, 1.243415e-05, -1.243415e-05, -1.02857e-05, 0, 0, 0,
  0, 0, 2.028637e-05, -4.036111e-05, -4.647492e-05, 4.647492e-05, 
    4.036111e-05, -2.028637e-05, 0, 0,
  0, -0.0001362561, -0.003977902, -0.002677063, -0.0008189927, 0.0008189927, 
    0.002677063, 0.003977902, 0.0001362561, 0,
  0.0002581271, -0.0009629345, -0.004511587, -0.002066068, -0.0003348062, 
    0.0003348062, 0.002066068, 0.004511587, 0.0009629345, -0.0002581271,
  0.0004235449, -0.001580223, -0.004630116, -0.000943519, -4.403178e-05, 
    4.403178e-05, 0.000943519, 0.004630116, 0.001580223, -0.0004235449,
  0.0004235449, -0.001580223, -0.004630116, -0.000943519, -4.403178e-05, 
    4.403178e-05, 0.000943519, 0.004630116, 0.001580223, -0.0004235449,
  0.0002581271, -0.0009629345, -0.004511587, -0.002066068, -0.0003348062, 
    0.0003348062, 0.002066068, 0.004511587, 0.0009629345, -0.0002581271,
  0, -0.0001362561, -0.003977902, -0.002677063, -0.0008189927, 0.0008189927, 
    0.002677063, 0.003977902, 0.0001362561, 0,
  0, 0, 2.028637e-05, -4.036111e-05, -4.647492e-05, 4.647492e-05, 
    4.036111e-05, -2.028637e-05, 0, 0,
  0, 0, 0, 1.02857e-05, 1.243415e-05, -1.243415e-05, -1.02857e-05, 0, 0, 0,
  0, 0, 0, 6.594866e-06, 8.130642e-06, -8.130642e-06, -6.594866e-06, 0, 0, 0,
  0, 0, 2.103172e-05, -2.552069e-05, -3.037642e-05, 3.037642e-05, 
    2.552069e-05, -2.103172e-05, 0, 0,
  0, -8.068501e-05, -0.002644493, -0.001780329, -0.0005451211, 0.0005451211, 
    0.001780329, 0.002644493, 8.068501e-05, 0,
  0.0001695268, -0.0006324865, -0.003004336, -0.001366226, -0.0002202333, 
    0.0002202333, 0.001366226, 0.003004336, 0.0006324865, -0.0001695268,
  0.0002789027, -0.00104065, -0.003085589, -0.0006189904, -2.871067e-05, 
    2.871067e-05, 0.0006189904, 0.003085589, 0.00104065, -0.0002789027,
  0.0002789027, -0.00104065, -0.003085589, -0.0006189904, -2.871067e-05, 
    2.871067e-05, 0.0006189904, 0.003085589, 0.00104065, -0.0002789027,
  0.0001695268, -0.0006324865, -0.003004336, -0.001366226, -0.0002202333, 
    0.0002202333, 0.001366226, 0.003004336, 0.0006324865, -0.0001695268,
  0, -8.068501e-05, -0.002644493, -0.001780329, -0.0005451211, 0.0005451211, 
    0.001780329, 0.002644493, 8.068501e-05, 0,
  0, 0, 2.103172e-05, -2.552069e-05, -3.037642e-05, 3.037642e-05, 
    2.552069e-05, -2.103172e-05, 0, 0,
  0, 0, 0, 6.594866e-06, 8.130642e-06, -8.130642e-06, -6.594866e-06, 0, 0, 0,
  0, 0, 0, 3.150988e-06, 3.961909e-06, -3.961909e-06, -3.150988e-06, 0, 0, 0,
  0, 0, 1.357571e-05, -1.200721e-05, -1.479293e-05, 1.479293e-05, 
    1.200721e-05, -1.357571e-05, 0, 0,
  0, -3.599225e-05, -0.001310641, -0.0008830633, -0.0002706518, 0.0002706518, 
    0.0008830633, 0.001310641, 3.599225e-05, 0,
  8.301486e-05, -0.0003097604, -0.001491929, -0.0006744439, -0.0001082485, 
    0.0001082485, 0.0006744439, 0.001491929, 0.0003097604, -8.301486e-05,
  0.0001368101, -0.0005105206, -0.001533798, -0.0003034991, -1.408372e-05, 
    1.408372e-05, 0.0003034991, 0.001533798, 0.0005105206, -0.0001368101,
  0.0001368101, -0.0005105206, -0.001533798, -0.0003034991, -1.408372e-05, 
    1.408372e-05, 0.0003034991, 0.001533798, 0.0005105206, -0.0001368101,
  8.301486e-05, -0.0003097604, -0.001491929, -0.0006744439, -0.0001082485, 
    0.0001082485, 0.0006744439, 0.001491929, 0.0003097604, -8.301486e-05,
  0, -3.599225e-05, -0.001310641, -0.0008830633, -0.0002706518, 0.0002706518, 
    0.0008830633, 0.001310641, 3.599225e-05, 0,
  0, 0, 1.357571e-05, -1.200721e-05, -1.479293e-05, 1.479293e-05, 
    1.200721e-05, -1.357571e-05, 0, 0,
  0, 0, 0, 3.150988e-06, 3.961909e-06, -3.961909e-06, -3.150988e-06, 0, 0, 0,
  0, 0, 0, 5.855569e-10, 3.119792e-10, -3.119792e-10, -5.855569e-10, 0, 0, 0,
  0, 0, -1.152815e-08, -4.240657e-09, -1.097102e-09, 1.097102e-09, 
    4.240657e-09, 1.152815e-08, 0, 0,
  0, -1.323016e-08, -2.346661e-08, -1.557423e-08, -4.872368e-09, 
    4.872368e-09, 1.557423e-08, 2.346661e-08, 1.323016e-08, 0,
  5.811907e-09, -2.378301e-08, -2.464363e-08, -1.542444e-08, -5.09584e-09, 
    5.09584e-09, 1.542444e-08, 2.464363e-08, 2.378301e-08, -5.811907e-09,
  7.001984e-09, -2.865949e-08, -2.544626e-08, -1.531423e-08, -5.821105e-09, 
    5.821105e-09, 1.531423e-08, 2.544626e-08, 2.865949e-08, -7.001984e-09,
  7.001984e-09, -2.865949e-08, -2.544626e-08, -1.531423e-08, -5.821105e-09, 
    5.821105e-09, 1.531423e-08, 2.544626e-08, 2.865949e-08, -7.001984e-09,
  5.811907e-09, -2.378301e-08, -2.464363e-08, -1.542444e-08, -5.09584e-09, 
    5.09584e-09, 1.542444e-08, 2.464363e-08, 2.378301e-08, -5.811907e-09,
  0, -1.323016e-08, -2.346661e-08, -1.557423e-08, -4.872368e-09, 
    4.872368e-09, 1.557423e-08, 2.346661e-08, 1.323016e-08, 0,
  0, 0, -1.152815e-08, -4.240657e-09, -1.097102e-09, 1.097102e-09, 
    4.240657e-09, 1.152815e-08, 0, 0,
  0, 0, 0, 5.855569e-10, 3.119792e-10, -3.119792e-10, -5.855569e-10, 0, 0, 0,
  0, 0, 0, 3.147144e-05, 2.767998e-05, -2.767998e-05, -3.147144e-05, 0, 0, 0,
  0, 0, -0.0002657369, -0.0001295755, -0.0001038073, 0.0001038073, 
    0.0001295755, 0.0002657369, 0, 0,
  0, -0.0007108127, -0.008294973, -0.005582972, -0.001717737, 0.001717737, 
    0.005582972, 0.008294973, 0.0007108127, 0,
  0.0006019049, -0.002244591, -0.009318897, -0.004578956, -0.0008463032, 
    0.0008463032, 0.004578956, 0.009318897, 0.002244591, -0.0006019049,
  0.0009306039, -0.003479775, -0.009625057, -0.002385959, -0.0001427074, 
    0.0001427074, 0.002385959, 0.009625057, 0.003479775, -0.0009306039,
  0.0009306039, -0.003479775, -0.009625057, -0.002385959, -0.0001427074, 
    0.0001427074, 0.002385959, 0.009625057, 0.003479775, -0.0009306039,
  0.0006019049, -0.002244591, -0.009318897, -0.004578956, -0.0008463032, 
    0.0008463032, 0.004578956, 0.009318897, 0.002244591, -0.0006019049,
  0, -0.0007108127, -0.008294973, -0.005582972, -0.001717737, 0.001717737, 
    0.005582972, 0.008294973, 0.0007108127, 0,
  0, 0, -0.0002657369, -0.0001295755, -0.0001038073, 0.0001038073, 
    0.0001295755, 0.0002657369, 0, 0,
  0, 0, 0, 3.147144e-05, 2.767998e-05, -2.767998e-05, -3.147144e-05, 0, 0, 0,
  0, 0, 0, 2.964231e-05, 2.744877e-05, -2.744877e-05, -2.964231e-05, 0, 0, 0,
  0, 0, -0.0002219629, -0.0001224955, -0.000102832, 0.000102832, 
    0.0001224955, 0.0002219629, 0, 0,
  0, -0.0006440201, -0.008224508, -0.005520921, -0.001694225, 0.001694225, 
    0.005520921, 0.008224508, 0.0006440201, 0,
  0.0005892332, -0.002197089, -0.009216779, -0.004501875, -0.0008165565, 
    0.0008165565, 0.004501875, 0.009216779, 0.002197089, -0.0005892332,
  0.0009190909, -0.00343237, -0.009496097, -0.0023104, -0.0001343212, 
    0.0001343212, 0.0023104, 0.009496097, 0.00343237, -0.0009190909,
  0.0009190909, -0.00343237, -0.009496097, -0.0023104, -0.0001343212, 
    0.0001343212, 0.0023104, 0.009496097, 0.00343237, -0.0009190909,
  0.0005892332, -0.002197089, -0.009216779, -0.004501875, -0.0008165565, 
    0.0008165565, 0.004501875, 0.009216779, 0.002197089, -0.0005892332,
  0, -0.0006440201, -0.008224508, -0.005520921, -0.001694225, 0.001694225, 
    0.005520921, 0.008224508, 0.0006440201, 0,
  0, 0, -0.0002219629, -0.0001224955, -0.000102832, 0.000102832, 
    0.0001224955, 0.0002219629, 0, 0,
  0, 0, 0, 2.964231e-05, 2.744877e-05, -2.744877e-05, -2.964231e-05, 0, 0, 0,
  0, 0, 0, 2.667872e-05, 2.664079e-05, -2.664079e-05, -2.667872e-05, 0, 0, 0,
  0, 0, -0.0001431774, -0.0001096674, -9.966083e-05, 9.966083e-05, 
    0.0001096674, 0.0001431774, 0, 0,
  0, -0.0005246762, -0.007956518, -0.005323435, -0.001625223, 0.001625223, 
    0.005323435, 0.007956518, 0.0005246762, 0,
  0.0005568951, -0.002076827, -0.008900011, -0.004267382, -0.0007479631, 
    0.0007479631, 0.004267382, 0.008900011, 0.002076827, -0.0005568951,
  0.0008832509, -0.003296289, -0.009123077, -0.002119857, -0.0001177278, 
    0.0001177278, 0.002119857, 0.009123077, 0.003296289, -0.0008832509,
  0.0008832509, -0.003296289, -0.009123077, -0.002119857, -0.0001177278, 
    0.0001177278, 0.002119857, 0.009123077, 0.003296289, -0.0008832509,
  0.0005568951, -0.002076827, -0.008900011, -0.004267382, -0.0007479631, 
    0.0007479631, 0.004267382, 0.008900011, 0.002076827, -0.0005568951,
  0, -0.0005246762, -0.007956518, -0.005323435, -0.001625223, 0.001625223, 
    0.005323435, 0.007956518, 0.0005246762, 0,
  0, 0, -0.0001431774, -0.0001096674, -9.966083e-05, 9.966083e-05, 
    0.0001096674, 0.0001431774, 0, 0,
  0, 0, 0, 2.667872e-05, 2.664079e-05, -2.664079e-05, -2.667872e-05, 0, 0, 0,
  0, 0, 0, 2.307964e-05, 2.435831e-05, -2.435831e-05, -2.307964e-05, 0, 0, 0,
  0, 0, -7.64058e-05, -9.385345e-05, -9.109949e-05, 9.109949e-05, 
    9.385345e-05, 7.64058e-05, 0, 0,
  0, -0.0004079585, -0.007352239, -0.004917953, -0.001498217, 0.001498217, 
    0.004917953, 0.007352239, 0.0004079585, 0,
  0.0005037647, -0.001878764, -0.008238082, -0.003885338, -0.00066039, 
    0.00066039, 0.003885338, 0.008238082, 0.001878764, -0.0005037647,
  0.0008088268, -0.00301774, -0.008422702, -0.001871772, -9.806082e-05, 
    9.806082e-05, 0.001871772, 0.008422702, 0.00301774, -0.0008088268,
  0.0008088268, -0.00301774, -0.008422702, -0.001871772, -9.806082e-05, 
    9.806082e-05, 0.001871772, 0.008422702, 0.00301774, -0.0008088268,
  0.0005037647, -0.001878764, -0.008238082, -0.003885338, -0.00066039, 
    0.00066039, 0.003885338, 0.008238082, 0.001878764, -0.0005037647,
  0, -0.0004079585, -0.007352239, -0.004917953, -0.001498217, 0.001498217, 
    0.004917953, 0.007352239, 0.0004079585, 0,
  0, 0, -7.64058e-05, -9.385345e-05, -9.109949e-05, 9.109949e-05, 
    9.385345e-05, 7.64058e-05, 0, 0,
  0, 0, 0, 2.307964e-05, 2.435831e-05, -2.435831e-05, -2.307964e-05, 0, 0, 0,
  0, 0, 0, 1.903953e-05, 2.092772e-05, -2.092772e-05, -1.903953e-05, 0, 0, 0,
  0, 0, -2.918386e-05, -7.647537e-05, -7.825991e-05, 7.825991e-05, 
    7.647537e-05, 2.918386e-05, 0, 0,
  0, -0.0003049664, -0.006424312, -0.004300881, -0.001310519, 0.001310519, 
    0.004300881, 0.006424312, 0.0003049664, 0,
  0.0004322374, -0.001612117, -0.007218394, -0.003362936, -0.0005603368, 
    0.0005603368, 0.003362936, 0.007218394, 0.001612117, -0.0004322374,
  0.0006996897, -0.002610353, -0.007378257, -0.001585539, -7.892161e-05, 
    7.892161e-05, 0.001585539, 0.007378257, 0.002610353, -0.0006996897,
  0.0006996897, -0.002610353, -0.007378257, -0.001585539, -7.892161e-05, 
    7.892161e-05, 0.001585539, 0.007378257, 0.002610353, -0.0006996897,
  0.0004322374, -0.001612117, -0.007218394, -0.003362936, -0.0005603368, 
    0.0005603368, 0.003362936, 0.007218394, 0.001612117, -0.0004322374,
  0, -0.0003049664, -0.006424312, -0.004300881, -0.001310519, 0.001310519, 
    0.004300881, 0.006424312, 0.0003049664, 0,
  0, 0, -2.918386e-05, -7.647537e-05, -7.825991e-05, 7.825991e-05, 
    7.647537e-05, 2.918386e-05, 0, 0,
  0, 0, 0, 1.903953e-05, 2.092772e-05, -2.092772e-05, -1.903953e-05, 0, 0, 0,
  0, 0, 0, 1.486524e-05, 1.686389e-05, -1.686389e-05, -1.486524e-05, 0, 0, 0,
  0, 0, 2.02782e-07, -5.895624e-05, -6.30493e-05, 6.30493e-05, 5.895624e-05, 
    -2.02782e-07, 0, 0,
  0, -0.0002173395, -0.005269258, -0.003530692, -0.00107686, 0.00107686, 
    0.003530692, 0.005269258, 0.0002173395, 0,
  0.0003490069, -0.001301814, -0.005936124, -0.002739154, -0.0004509174, 
    0.0004509174, 0.002739154, 0.005936124, 0.001301814, -0.0003490069,
  0.0005682205, -0.002119897, -0.00607133, -0.001272735, -6.133533e-05, 
    6.133533e-05, 0.001272735, 0.00607133, 0.002119897, -0.0005682205,
  0.0005682205, -0.002119897, -0.00607133, -0.001272735, -6.133533e-05, 
    6.133533e-05, 0.001272735, 0.00607133, 0.002119897, -0.0005682205,
  0.0003490069, -0.001301814, -0.005936124, -0.002739154, -0.0004509174, 
    0.0004509174, 0.002739154, 0.005936124, 0.001301814, -0.0003490069,
  0, -0.0002173395, -0.005269258, -0.003530692, -0.00107686, 0.00107686, 
    0.003530692, 0.005269258, 0.0002173395, 0,
  0, 0, 2.02782e-07, -5.895624e-05, -6.30493e-05, 6.30493e-05, 5.895624e-05, 
    -2.02782e-07, 0, 0,
  0, 0, 0, 1.486524e-05, 1.686389e-05, -1.686389e-05, -1.486524e-05, 0, 0, 0,
  0, 0, 0, 1.078954e-05, 1.253975e-05, -1.253975e-05, -1.078954e-05, 0, 0, 0,
  0, 0, 1.449837e-05, -4.224362e-05, -4.68675e-05, 4.68675e-05, 4.224362e-05, 
    -1.449837e-05, 0, 0,
  0, -0.0001452263, -0.003986346, -0.00267257, -0.0008159337, 0.0008159337, 
    0.00267257, 0.003986346, 0.0001452263, 0,
  0.000260449, -0.0009715913, -0.004500266, -0.00205993, -0.0003365328, 
    0.0003365328, 0.00205993, 0.004500266, 0.0009715913, -0.000260449,
  0.0004257144, -0.001588321, -0.004606354, -0.0009472928, -4.491138e-05, 
    4.491138e-05, 0.0009472928, 0.004606354, 0.001588321, -0.0004257144,
  0.0004257144, -0.001588321, -0.004606354, -0.0009472928, -4.491138e-05, 
    4.491138e-05, 0.0009472928, 0.004606354, 0.001588321, -0.0004257144,
  0.000260449, -0.0009715913, -0.004500266, -0.00205993, -0.0003365328, 
    0.0003365328, 0.00205993, 0.004500266, 0.0009715913, -0.000260449,
  0, -0.0001452263, -0.003986346, -0.00267257, -0.0008159337, 0.0008159337, 
    0.00267257, 0.003986346, 0.0001452263, 0,
  0, 0, 1.449837e-05, -4.224362e-05, -4.68675e-05, 4.68675e-05, 4.224362e-05, 
    -1.449837e-05, 0, 0,
  0, 0, 0, 1.078954e-05, 1.253975e-05, -1.253975e-05, -1.078954e-05, 0, 0, 0,
  0, 0, 0, 6.926054e-06, 8.20167e-06, -8.20167e-06, -6.926054e-06, 0, 0, 0,
  0, 0, 1.717206e-05, -2.675768e-05, -3.064086e-05, 3.064086e-05, 
    2.675768e-05, -1.717206e-05, 0, 0,
  0, -8.680863e-05, -0.002652172, -0.001778646, -0.0005434534, 0.0005434534, 
    0.001778646, 0.002652172, 8.680863e-05, 0,
  0.0001711433, -0.0006385141, -0.002999044, -0.001362896, -0.0002215119, 
    0.0002215119, 0.001362896, 0.002999044, 0.0006385141, -0.0001711433,
  0.0002804244, -0.001046328, -0.003071944, -0.0006218205, -2.930621e-05, 
    2.930621e-05, 0.0006218205, 0.003071944, 0.001046328, -0.0002804244,
  0.0002804244, -0.001046328, -0.003071944, -0.0006218205, -2.930621e-05, 
    2.930621e-05, 0.0006218205, 0.003071944, 0.001046328, -0.0002804244,
  0.0001711433, -0.0006385141, -0.002999044, -0.001362896, -0.0002215119, 
    0.0002215119, 0.001362896, 0.002999044, 0.0006385141, -0.0001711433,
  0, -8.680863e-05, -0.002652172, -0.001778646, -0.0005434534, 0.0005434534, 
    0.001778646, 0.002652172, 8.680863e-05, 0,
  0, 0, 1.717206e-05, -2.675768e-05, -3.064086e-05, 3.064086e-05, 
    2.675768e-05, -1.717206e-05, 0, 0,
  0, 0, 0, 6.926054e-06, 8.20167e-06, -8.20167e-06, -6.926054e-06, 0, 0, 0,
  0, 0, 0, 3.30618e-06, 3.997906e-06, -3.997906e-06, -3.30618e-06, 0, 0, 0,
  0, 0, 1.176195e-05, -1.258667e-05, -1.492714e-05, 1.492714e-05, 
    1.258667e-05, -1.176195e-05, 0, 0,
  0, -3.896345e-05, -0.001315608, -0.0008832358, -0.0002701678, 0.0002701678, 
    0.0008832358, 0.001315608, 3.896345e-05, 0,
  8.384304e-05, -0.0003128497, -0.001491015, -0.000673676, -0.0001090037, 
    0.0001090037, 0.000673676, 0.001491015, 0.0003128497, -8.384304e-05,
  0.0001376203, -0.0005135435, -0.001528998, -0.0003052508, -1.43951e-05, 
    1.43951e-05, 0.0003052508, 0.001528998, 0.0005135435, -0.0001376203,
  0.0001376203, -0.0005135435, -0.001528998, -0.0003052508, -1.43951e-05, 
    1.43951e-05, 0.0003052508, 0.001528998, 0.0005135435, -0.0001376203,
  8.384304e-05, -0.0003128497, -0.001491015, -0.000673676, -0.0001090037, 
    0.0001090037, 0.000673676, 0.001491015, 0.0003128497, -8.384304e-05,
  0, -3.896345e-05, -0.001315608, -0.0008832358, -0.0002701678, 0.0002701678, 
    0.0008832358, 0.001315608, 3.896345e-05, 0,
  0, 0, 1.176195e-05, -1.258667e-05, -1.492714e-05, 1.492714e-05, 
    1.258667e-05, -1.176195e-05, 0, 0,
  0, 0, 0, 3.30618e-06, 3.997906e-06, -3.997906e-06, -3.30618e-06, 0, 0, 0,
  0, 0, 0, 5.857667e-10, 3.120892e-10, -3.120892e-10, -5.857667e-10, 0, 0, 0,
  0, 0, -1.15415e-08, -4.246539e-09, -1.097673e-09, 1.097673e-09, 
    4.246539e-09, 1.15415e-08, 0, 0,
  0, -1.32585e-08, -2.346004e-08, -1.556134e-08, -4.869617e-09, 4.869617e-09, 
    1.556134e-08, 2.346004e-08, 1.32585e-08, 0,
  5.815344e-09, -2.381267e-08, -2.459297e-08, -1.540685e-08, -5.098232e-09, 
    5.098232e-09, 1.540685e-08, 2.459297e-08, 2.381267e-08, -5.815344e-09,
  7.002647e-09, -2.868336e-08, -2.537498e-08, -1.532166e-08, -5.842038e-09, 
    5.842038e-09, 1.532166e-08, 2.537498e-08, 2.868336e-08, -7.002647e-09,
  7.002647e-09, -2.868336e-08, -2.537498e-08, -1.532166e-08, -5.842038e-09, 
    5.842038e-09, 1.532166e-08, 2.537498e-08, 2.868336e-08, -7.002647e-09,
  5.815344e-09, -2.381267e-08, -2.459297e-08, -1.540685e-08, -5.098232e-09, 
    5.098232e-09, 1.540685e-08, 2.459297e-08, 2.381267e-08, -5.815344e-09,
  0, -1.32585e-08, -2.346004e-08, -1.556134e-08, -4.869617e-09, 4.869617e-09, 
    1.556134e-08, 2.346004e-08, 1.32585e-08, 0,
  0, 0, -1.15415e-08, -4.246539e-09, -1.097673e-09, 1.097673e-09, 
    4.246539e-09, 1.15415e-08, 0, 0,
  0, 0, 0, 5.857667e-10, 3.120892e-10, -3.120892e-10, -5.857667e-10, 0, 0, 0,
  0, 0, 0, 3.247311e-05, 2.790047e-05, -2.790047e-05, -3.247311e-05, 0, 0, 0,
  0, 0, -0.0002768362, -0.0001333559, -0.0001046175, 0.0001046175, 
    0.0001333559, 0.0002768362, 0, 0,
  0, -0.00072758, -0.008301422, -0.005568251, -0.001709754, 0.001709754, 
    0.005568251, 0.008301422, 0.00072758, 0,
  0.0006061294, -0.002260444, -0.009286314, -0.004563344, -0.0008484946, 
    0.0008484946, 0.004563344, 0.009286314, 0.002260444, -0.0006061294,
  0.0009345636, -0.00349472, -0.009566539, -0.002390856, -0.000145277, 
    0.000145277, 0.002390856, 0.009566539, 0.00349472, -0.0009345636,
  0.0009345636, -0.00349472, -0.009566539, -0.002390856, -0.000145277, 
    0.000145277, 0.002390856, 0.009566539, 0.00349472, -0.0009345636,
  0.0006061294, -0.002260444, -0.009286314, -0.004563344, -0.0008484946, 
    0.0008484946, 0.004563344, 0.009286314, 0.002260444, -0.0006061294,
  0, -0.00072758, -0.008301422, -0.005568251, -0.001709754, 0.001709754, 
    0.005568251, 0.008301422, 0.00072758, 0,
  0, 0, -0.0002768362, -0.0001333559, -0.0001046175, 0.0001046175, 
    0.0001333559, 0.0002768362, 0, 0,
  0, 0, 0, 3.247311e-05, 2.790047e-05, -2.790047e-05, -3.247311e-05, 0, 0, 0,
  0, 0, 0, 3.064858e-05, 2.766737e-05, -2.766737e-05, -3.064858e-05, 0, 0, 0,
  0, 0, -0.0002331512, -0.0001262809, -0.0001036354, 0.0001036354, 
    0.0001262809, 0.0002331512, 0, 0,
  0, -0.0006609037, -0.008230937, -0.005506466, -0.001686466, 0.001686466, 
    0.005506466, 0.008230937, 0.0006609037, 0,
  0.0005934635, -0.002212907, -0.009184726, -0.004486478, -0.0008188451, 
    0.0008188451, 0.004486478, 0.009184726, 0.002212907, -0.0005934635,
  0.000923071, -0.003447313, -0.009438962, -0.002315367, -0.0001367709, 
    0.0001367709, 0.002315367, 0.009438962, 0.003447313, -0.000923071,
  0.000923071, -0.003447313, -0.009438962, -0.002315367, -0.0001367709, 
    0.0001367709, 0.002315367, 0.009438962, 0.003447313, -0.000923071,
  0.0005934635, -0.002212907, -0.009184726, -0.004486478, -0.0008188451, 
    0.0008188451, 0.004486478, 0.009184726, 0.002212907, -0.0005934635,
  0, -0.0006609037, -0.008230937, -0.005506466, -0.001686466, 0.001686466, 
    0.005506466, 0.008230937, 0.0006609037, 0,
  0, 0, -0.0002331512, -0.0001262809, -0.0001036354, 0.0001036354, 
    0.0001262809, 0.0002331512, 0, 0,
  0, 0, 0, 3.064858e-05, 2.766737e-05, -2.766737e-05, -3.064858e-05, 0, 0, 0,
  0, 0, 0, 2.767257e-05, 2.685105e-05, -2.685105e-05, -2.767257e-05, 0, 0, 0,
  0, 0, -0.0001542188, -0.0001133935, -0.0001004356, 0.0001004356, 
    0.0001133935, 0.0001542188, 0, 0,
  0, -0.0005412701, -0.007963161, -0.005309715, -0.001617949, 0.001617949, 
    0.005309715, 0.007963161, 0.0005412701, 0,
  0.0005610802, -0.002092445, -0.008869411, -0.004252854, -0.0007504071, 
    0.0007504071, 0.004252854, 0.008869411, 0.002092445, -0.0005610802,
  0.0008871742, -0.003310974, -0.009069029, -0.002125125, -0.0001198822, 
    0.0001198822, 0.002125125, 0.009069029, 0.003310974, -0.0008871742,
  0.0008871742, -0.003310974, -0.009069029, -0.002125125, -0.0001198822, 
    0.0001198822, 0.002125125, 0.009069029, 0.003310974, -0.0008871742,
  0.0005610802, -0.002092445, -0.008869411, -0.004252854, -0.0007504071, 
    0.0007504071, 0.004252854, 0.008869411, 0.002092445, -0.0005610802,
  0, -0.0005412701, -0.007963161, -0.005309715, -0.001617949, 0.001617949, 
    0.005309715, 0.007963161, 0.0005412701, 0,
  0, 0, -0.0001542188, -0.0001133935, -0.0001004356, 0.0001004356, 
    0.0001133935, 0.0001542188, 0, 0,
  0, 0, 0, 2.767257e-05, 2.685105e-05, -2.685105e-05, -2.767257e-05, 0, 0, 0,
  0, 0, 0, 2.400551e-05, 2.455148e-05, -2.455148e-05, -2.400551e-05, 0, 0, 0,
  0, 0, -8.674272e-05, -9.731921e-05, -9.181334e-05, 9.181334e-05, 
    9.731921e-05, 8.674272e-05, 0, 0,
  0, -0.0004234944, -0.007359335, -0.004905664, -0.001491658, 0.001491658, 
    0.004905664, 0.007359335, 0.0004234944, 0,
  0.000507704, -0.001893454, -0.008210418, -0.003872271, -0.0006628838, 
    0.0006628838, 0.003872271, 0.008210418, 0.001893454, -0.000507704,
  0.0008125075, -0.003031498, -0.008373619, -0.001877165, -9.98738e-05, 
    9.98738e-05, 0.001877165, 0.008373619, 0.003031498, -0.0008125075,
  0.0008125075, -0.003031498, -0.008373619, -0.001877165, -9.98738e-05, 
    9.98738e-05, 0.001877165, 0.008373619, 0.003031498, -0.0008125075,
  0.000507704, -0.001893454, -0.008210418, -0.003872271, -0.0006628838, 
    0.0006628838, 0.003872271, 0.008210418, 0.001893454, -0.000507704,
  0, -0.0004234944, -0.007359335, -0.004905664, -0.001491658, 0.001491658, 
    0.004905664, 0.007359335, 0.0004234944, 0,
  0, 0, -8.674272e-05, -9.731921e-05, -9.181334e-05, 9.181334e-05, 
    9.731921e-05, 8.674272e-05, 0, 0,
  0, 0, 0, 2.400551e-05, 2.455148e-05, -2.455148e-05, -2.400551e-05, 0, 0, 0,
  0, 0, 0, 1.984986e-05, 2.109633e-05, -2.109633e-05, -1.984986e-05, 0, 0, 0,
  0, 0, -3.829163e-05, -7.950608e-05, -7.888443e-05, 7.888443e-05, 
    7.950608e-05, 3.829163e-05, 0, 0,
  0, -0.0003187215, -0.006431939, -0.004290752, -0.001304943, 0.001304943, 
    0.004290752, 0.006431939, 0.0003187215, 0,
  0.0004357429, -0.001625186, -0.007195233, -0.003351852, -0.000562699, 
    0.000562699, 0.003351852, 0.007195233, 0.001625186, -0.0004357429,
  0.0007029631, -0.002622579, -0.007336242, -0.001590661, -8.040916e-05, 
    8.040916e-05, 0.001590661, 0.007336242, 0.002622579, -0.0007029631,
  0.0007029631, -0.002622579, -0.007336242, -0.001590661, -8.040916e-05, 
    8.040916e-05, 0.001590661, 0.007336242, 0.002622579, -0.0007029631,
  0.0004357429, -0.001625186, -0.007195233, -0.003351852, -0.000562699, 
    0.000562699, 0.003351852, 0.007195233, 0.001625186, -0.0004357429,
  0, -0.0003187215, -0.006431939, -0.004290752, -0.001304943, 0.001304943, 
    0.004290752, 0.006431939, 0.0003187215, 0,
  0, 0, -3.829163e-05, -7.950608e-05, -7.888443e-05, 7.888443e-05, 
    7.950608e-05, 3.829163e-05, 0, 0,
  0, 0, 0, 1.984986e-05, 2.109633e-05, -2.109633e-05, -1.984986e-05, 0, 0, 0,
  0, 0, 0, 1.552998e-05, 1.700224e-05, -1.700224e-05, -1.552998e-05, 0, 0, 0,
  0, 0, -7.34213e-06, -6.144099e-05, -6.356273e-05, 6.356273e-05, 
    6.144099e-05, 7.34213e-06, 0, 0,
  0, -0.0002288451, -0.005277331, -0.003523243, -0.001072489, 0.001072489, 
    0.003523243, 0.005277331, 0.0002288451, 0,
  0.0003519526, -0.001312796, -0.005918587, -0.00273045, -0.0004529995, 
    0.0004529995, 0.00273045, 0.005918587, 0.001312796, -0.0003519526,
  0.000570968, -0.002130154, -0.006038046, -0.001277258, -6.251538e-05, 
    6.251538e-05, 0.001277258, 0.006038046, 0.002130154, -0.000570968,
  0.000570968, -0.002130154, -0.006038046, -0.001277258, -6.251538e-05, 
    6.251538e-05, 0.001277258, 0.006038046, 0.002130154, -0.000570968,
  0.0003519526, -0.001312796, -0.005918587, -0.00273045, -0.0004529995, 
    0.0004529995, 0.00273045, 0.005918587, 0.001312796, -0.0003519526,
  0, -0.0002288451, -0.005277331, -0.003523243, -0.001072489, 0.001072489, 
    0.003523243, 0.005277331, 0.0002288451, 0,
  0, 0, -7.34213e-06, -6.144099e-05, -6.356273e-05, 6.356273e-05, 
    6.144099e-05, 7.34213e-06, 0, 0,
  0, 0, 0, 1.552998e-05, 1.700224e-05, -1.700224e-05, -1.552998e-05, 0, 0, 0,
  0, 0, 0, 1.129161e-05, 1.264471e-05, -1.264471e-05, -1.129161e-05, 0, 0, 0,
  0, 0, 8.722372e-06, -4.411942e-05, -4.725766e-05, 4.725766e-05, 
    4.411942e-05, -8.722372e-06, 0, 0,
  0, -0.0001541701, -0.003994514, -0.002668035, -0.0008129022, 0.0008129022, 
    0.002668035, 0.003994514, 0.0001541701, 0,
  0.0002627548, -0.0009801878, -0.004488886, -0.002053865, -0.0003382375, 
    0.0003382375, 0.002053865, 0.004488886, 0.0009801878, -0.0002627548,
  0.0004278635, -0.001596342, -0.004582806, -0.0009510084, -4.579626e-05, 
    4.579626e-05, 0.0009510084, 0.004582806, 0.001596342, -0.0004278635,
  0.0004278635, -0.001596342, -0.004582806, -0.0009510084, -4.579626e-05, 
    4.579626e-05, 0.0009510084, 0.004582806, 0.001596342, -0.0004278635,
  0.0002627548, -0.0009801878, -0.004488886, -0.002053865, -0.0003382375, 
    0.0003382375, 0.002053865, 0.004488886, 0.0009801878, -0.0002627548,
  0, -0.0001541701, -0.003994514, -0.002668035, -0.0008129022, 0.0008129022, 
    0.002668035, 0.003994514, 0.0001541701, 0,
  0, 0, 8.722372e-06, -4.411942e-05, -4.725766e-05, 4.725766e-05, 
    4.411942e-05, -8.722372e-06, 0, 0,
  0, 0, 0, 1.129161e-05, 1.264471e-05, -1.264471e-05, -1.129161e-05, 0, 0, 0,
  0, 0, 0, 7.255041e-06, 8.272434e-06, -8.272434e-06, -7.255041e-06, 0, 0, 0,
  0, 0, 1.334456e-05, -2.798641e-05, -3.090431e-05, 3.090431e-05, 
    2.798641e-05, -1.334456e-05, 0, 0,
  0, -9.286299e-05, -0.002659449, -0.001776851, -0.0005417906, 0.0005417906, 
    0.001776851, 0.002659449, 9.286299e-05, 0,
  0.0001727396, -0.0006444664, -0.002993557, -0.001359622, -0.000222772, 
    0.000222772, 0.001359622, 0.002993557, 0.0006444664, -0.0001727396,
  0.0002819296, -0.001051945, -0.003058342, -0.0006246124, -2.990525e-05, 
    2.990525e-05, 0.0006246124, 0.003058342, 0.001051945, -0.0002819296,
  0.0002819296, -0.001051945, -0.003058342, -0.0006246124, -2.990525e-05, 
    2.990525e-05, 0.0006246124, 0.003058342, 0.001051945, -0.0002819296,
  0.0001727396, -0.0006444664, -0.002993557, -0.001359622, -0.000222772, 
    0.000222772, 0.001359622, 0.002993557, 0.0006444664, -0.0001727396,
  0, -9.286299e-05, -0.002659449, -0.001776851, -0.0005417906, 0.0005417906, 
    0.001776851, 0.002659449, 9.286299e-05, 0,
  0, 0, 1.334456e-05, -2.798641e-05, -3.090431e-05, 3.090431e-05, 
    2.798641e-05, -1.334456e-05, 0, 0,
  0, 0, 0, 7.255041e-06, 8.272434e-06, -8.272434e-06, -7.255041e-06, 0, 0, 0,
  0, 0, 0, 3.460302e-06, 4.033622e-06, -4.033622e-06, -3.460302e-06, 0, 0, 0,
  0, 0, 9.967926e-06, -1.316213e-05, -1.50603e-05, 1.50603e-05, 1.316213e-05, 
    -9.967926e-06, 0, 0,
  0, -4.188015e-05, -0.00132016, -0.0008832128, -0.0002696476, 0.0002696476, 
    0.0008832128, 0.00132016, 4.188015e-05, 0,
  8.465277e-05, -0.0003158701, -0.001489761, -0.000672873, -0.0001097427, 
    0.0001097427, 0.000672873, 0.001489761, 0.0003158701, -8.465277e-05,
  0.000138414, -0.0005165051, -0.001523985, -0.0003069691, -1.470675e-05, 
    1.470675e-05, 0.0003069691, 0.001523985, 0.0005165051, -0.000138414,
  0.000138414, -0.0005165051, -0.001523985, -0.0003069691, -1.470675e-05, 
    1.470675e-05, 0.0003069691, 0.001523985, 0.0005165051, -0.000138414,
  8.465277e-05, -0.0003158701, -0.001489761, -0.000672873, -0.0001097427, 
    0.0001097427, 0.000672873, 0.001489761, 0.0003158701, -8.465277e-05,
  0, -4.188015e-05, -0.00132016, -0.0008832128, -0.0002696476, 0.0002696476, 
    0.0008832128, 0.00132016, 4.188015e-05, 0,
  0, 0, 9.967926e-06, -1.316213e-05, -1.50603e-05, 1.50603e-05, 1.316213e-05, 
    -9.967926e-06, 0, 0,
  0, 0, 0, 3.460302e-06, 4.033622e-06, -4.033622e-06, -3.460302e-06, 0, 0, 0,
  0, 0, 0, 5.859639e-10, 3.12195e-10, -3.12195e-10, -5.859639e-10, 0, 0, 0,
  0, 0, -1.155473e-08, -4.252366e-09, -1.098231e-09, 1.098231e-09, 
    4.252366e-09, 1.155473e-08, 0, 0,
  0, -1.328672e-08, -2.345341e-08, -1.554851e-08, -4.866877e-09, 
    4.866877e-09, 1.554851e-08, 2.345341e-08, 1.328672e-08, 0,
  5.818711e-09, -2.384211e-08, -2.454256e-08, -1.538936e-08, -5.100642e-09, 
    5.100642e-09, 1.538936e-08, 2.454256e-08, 2.384211e-08, -5.818711e-09,
  7.003219e-09, -2.870693e-08, -2.530428e-08, -1.532886e-08, -5.862804e-09, 
    5.862804e-09, 1.532886e-08, 2.530428e-08, 2.870693e-08, -7.003219e-09,
  7.003219e-09, -2.870693e-08, -2.530428e-08, -1.532886e-08, -5.862804e-09, 
    5.862804e-09, 1.532886e-08, 2.530428e-08, 2.870693e-08, -7.003219e-09,
  5.818711e-09, -2.384211e-08, -2.454256e-08, -1.538936e-08, -5.100642e-09, 
    5.100642e-09, 1.538936e-08, 2.454256e-08, 2.384211e-08, -5.818711e-09,
  0, -1.328672e-08, -2.345341e-08, -1.554851e-08, -4.866877e-09, 
    4.866877e-09, 1.554851e-08, 2.345341e-08, 1.328672e-08, 0,
  0, 0, -1.155473e-08, -4.252366e-09, -1.098231e-09, 1.098231e-09, 
    4.252366e-09, 1.155473e-08, 0, 0,
  0, 0, 0, 5.859639e-10, 3.12195e-10, -3.12195e-10, -5.859639e-10, 0, 0, 0,
  0, 0, 0, 3.347251e-05, 2.81193e-05, -2.81193e-05, -3.347251e-05, 0, 0, 0,
  0, 0, -0.0002879208, -0.0001371278, -0.0001054216, 0.0001054216, 
    0.0001371278, 0.0002879208, 0, 0,
  0, -0.0007443273, -0.008307651, -0.005553571, -0.001701849, 0.001701849, 
    0.005553571, 0.008307651, 0.0007443273, 0,
  0.0006103343, -0.002276226, -0.00925385, -0.004547864, -0.0008506518, 
    0.0008506518, 0.004547864, 0.00925385, 0.002276226, -0.0006103343,
  0.0009384871, -0.003509531, -0.009508641, -0.002395635, -0.0001478502, 
    0.0001478502, 0.002395635, 0.009508641, 0.003509531, -0.0009384871,
  0.0009384871, -0.003509531, -0.009508641, -0.002395635, -0.0001478502, 
    0.0001478502, 0.002395635, 0.009508641, 0.003509531, -0.0009384871,
  0.0006103343, -0.002276226, -0.00925385, -0.004547864, -0.0008506518, 
    0.0008506518, 0.004547864, 0.00925385, 0.002276226, -0.0006103343,
  0, -0.0007443273, -0.008307651, -0.005553571, -0.001701849, 0.001701849, 
    0.005553571, 0.008307651, 0.0007443273, 0,
  0, 0, -0.0002879208, -0.0001371278, -0.0001054216, 0.0001054216, 
    0.0001371278, 0.0002879208, 0, 0,
  0, 0, 0, 3.347251e-05, 2.81193e-05, -2.81193e-05, -3.347251e-05, 0, 0, 0,
  0, 0, 0, 3.165267e-05, 2.788437e-05, -2.788437e-05, -3.165267e-05, 0, 0, 0,
  0, 0, -0.0002443254, -0.000130058, -0.0001044329, 0.0001044329, 
    0.000130058, 0.0002443254, 0, 0,
  0, -0.0006777684, -0.008237146, -0.00549205, -0.001678783, 0.001678783, 
    0.00549205, 0.008237146, 0.0006777684, 0,
  0.0005976752, -0.002228657, -0.009152789, -0.004471213, -0.000821099, 
    0.000821099, 0.004471213, 0.009152789, 0.002228657, -0.0005976752,
  0.0009270158, -0.003462126, -0.00938243, -0.002320217, -0.0001392249, 
    0.0001392249, 0.002320217, 0.00938243, 0.003462126, -0.0009270158,
  0.0009270158, -0.003462126, -0.00938243, -0.002320217, -0.0001392249, 
    0.0001392249, 0.002320217, 0.00938243, 0.003462126, -0.0009270158,
  0.0005976752, -0.002228657, -0.009152789, -0.004471213, -0.000821099, 
    0.000821099, 0.004471213, 0.009152789, 0.002228657, -0.0005976752,
  0, -0.0006777684, -0.008237146, -0.00549205, -0.001678783, 0.001678783, 
    0.00549205, 0.008237146, 0.0006777684, 0,
  0, 0, -0.0002443254, -0.000130058, -0.0001044329, 0.0001044329, 
    0.000130058, 0.0002443254, 0, 0,
  0, 0, 0, 3.165267e-05, 2.788437e-05, -2.788437e-05, -3.165267e-05, 0, 0, 0,
  0, 0, 0, 2.866435e-05, 2.705974e-05, -2.705974e-05, -2.866435e-05, 0, 0, 0,
  0, 0, -0.0001652497, -0.0001171117, -0.0001012046, 0.0001012046, 
    0.0001171117, 0.0001652497, 0, 0,
  0, -0.0005578496, -0.007969586, -0.005296031, -0.001610746, 0.001610746, 
    0.005296031, 0.007969586, 0.0005578496, 0,
  0.0005652474, -0.002107996, -0.008838919, -0.004238452, -0.0007528162, 
    0.0007528162, 0.004238452, 0.008838919, 0.002107996, -0.0005652474,
  0.000891063, -0.003325532, -0.009015546, -0.00213028, -0.0001220418, 
    0.0001220418, 0.00213028, 0.009015546, 0.003325532, -0.000891063,
  0.000891063, -0.003325532, -0.009015546, -0.00213028, -0.0001220418, 
    0.0001220418, 0.00213028, 0.009015546, 0.003325532, -0.000891063,
  0.0005652474, -0.002107996, -0.008838919, -0.004238452, -0.0007528162, 
    0.0007528162, 0.004238452, 0.008838919, 0.002107996, -0.0005652474,
  0, -0.0005578496, -0.007969586, -0.005296031, -0.001610746, 0.001610746, 
    0.005296031, 0.007969586, 0.0005578496, 0,
  0, 0, -0.0001652497, -0.0001171117, -0.0001012046, 0.0001012046, 
    0.0001171117, 0.0001652497, 0, 0,
  0, 0, 0, 2.866435e-05, 2.705974e-05, -2.705974e-05, -2.866435e-05, 0, 0, 0,
  0, 0, 0, 2.492957e-05, 2.474323e-05, -2.474323e-05, -2.492957e-05, 0, 0, 0,
  0, 0, -9.707255e-05, -0.000100778, -9.252194e-05, 9.252194e-05, 
    0.000100778, 9.707255e-05, 0, 0,
  0, -0.0004390201, -0.007366215, -0.004893403, -0.001485162, 0.001485162, 
    0.004893403, 0.007366215, 0.0004390201, 0,
  0.0005116269, -0.001908083, -0.00818284, -0.003859318, -0.0006653439, 
    0.0006653439, 0.003859318, 0.00818284, 0.001908083, -0.0005116269,
  0.0008161564, -0.003045139, -0.008325042, -0.001882452, -0.0001016929, 
    0.0001016929, 0.001882452, 0.008325042, 0.003045139, -0.0008161564,
  0.0008161564, -0.003045139, -0.008325042, -0.001882452, -0.0001016929, 
    0.0001016929, 0.001882452, 0.008325042, 0.003045139, -0.0008161564,
  0.0005116269, -0.001908083, -0.00818284, -0.003859318, -0.0006653439, 
    0.0006653439, 0.003859318, 0.00818284, 0.001908083, -0.0005116269,
  0, -0.0004390201, -0.007366215, -0.004893403, -0.001485162, 0.001485162, 
    0.004893403, 0.007366215, 0.0004390201, 0,
  0, 0, -9.707255e-05, -0.000100778, -9.252194e-05, 9.252194e-05, 
    0.000100778, 9.707255e-05, 0, 0,
  0, 0, 0, 2.492957e-05, 2.474323e-05, -2.474323e-05, -2.492957e-05, 0, 0, 0,
  0, 0, 0, 2.065873e-05, 2.126374e-05, -2.126374e-05, -2.065873e-05, 0, 0, 0,
  0, 0, -4.739587e-05, -8.253117e-05, -7.950452e-05, 7.950452e-05, 
    8.253117e-05, 4.739587e-05, 0, 0,
  0, -0.00033247, -0.006439356, -0.004280637, -0.001299421, 0.001299421, 
    0.004280637, 0.006439356, 0.00033247, 0,
  0.0004392341, -0.001638202, -0.007172128, -0.003340868, -0.0005650306, 
    0.0005650306, 0.003340868, 0.007172128, 0.001638202, -0.0004392341,
  0.0007062089, -0.002634703, -0.007294649, -0.001595689, -8.190312e-05, 
    8.190312e-05, 0.001595689, 0.007294649, 0.002634703, -0.0007062089,
  0.0007062089, -0.002634703, -0.007294649, -0.001595689, -8.190312e-05, 
    8.190312e-05, 0.001595689, 0.007294649, 0.002634703, -0.0007062089,
  0.0004392341, -0.001638202, -0.007172128, -0.003340868, -0.0005650306, 
    0.0005650306, 0.003340868, 0.007172128, 0.001638202, -0.0004392341,
  0, -0.00033247, -0.006439356, -0.004280637, -0.001299421, 0.001299421, 
    0.004280637, 0.006439356, 0.00033247, 0,
  0, 0, -4.739587e-05, -8.253117e-05, -7.950452e-05, 7.950452e-05, 
    8.253117e-05, 4.739587e-05, 0, 0,
  0, 0, 0, 2.065873e-05, 2.126374e-05, -2.126374e-05, -2.065873e-05, 0, 0, 0,
  0, 0, 0, 1.619353e-05, 1.713968e-05, -1.713968e-05, -1.619353e-05, 0, 0, 0,
  0, 0, -1.488402e-05, -6.392113e-05, -6.40728e-05, 6.40728e-05, 
    6.392113e-05, 1.488402e-05, 0, 0,
  0, -0.0002403419, -0.00528519, -0.003515788, -0.001068158, 0.001068158, 
    0.003515788, 0.00528519, 0.0002403419, 0,
  0.000354886, -0.001323731, -0.005901063, -0.002721828, -0.0004550555, 
    0.0004550555, 0.002721828, 0.005901063, 0.001323731, -0.000354886,
  0.0005736933, -0.002140329, -0.006005088, -0.001281703, -6.370142e-05, 
    6.370142e-05, 0.001281703, 0.006005088, 0.002140329, -0.0005736933,
  0.0005736933, -0.002140329, -0.006005088, -0.001281703, -6.370142e-05, 
    6.370142e-05, 0.001281703, 0.006005088, 0.002140329, -0.0005736933,
  0.000354886, -0.001323731, -0.005901063, -0.002721828, -0.0004550555, 
    0.0004550555, 0.002721828, 0.005901063, 0.001323731, -0.000354886,
  0, -0.0002403419, -0.00528519, -0.003515788, -0.001068158, 0.001068158, 
    0.003515788, 0.00528519, 0.0002403419, 0,
  0, 0, -1.488402e-05, -6.392113e-05, -6.40728e-05, 6.40728e-05, 
    6.392113e-05, 1.488402e-05, 0, 0,
  0, 0, 0, 1.619353e-05, 1.713968e-05, -1.713968e-05, -1.619353e-05, 0, 0, 0,
  0, 0, 0, 1.179233e-05, 1.274914e-05, -1.274914e-05, -1.179233e-05, 0, 0, 0,
  0, 0, 2.959485e-06, -4.599014e-05, -4.764587e-05, 4.764587e-05, 
    4.599014e-05, -2.959485e-06, 0, 0,
  0, -0.0001630833, -0.004002416, -0.002663461, -0.0008098975, 0.0008098975, 
    0.002663461, 0.004002416, 0.0001630833, 0,
  0.0002650476, -0.0009887358, -0.004477448, -0.002047871, -0.0003399205, 
    0.0003399205, 0.002047871, 0.004477448, 0.0009887358, -0.0002650476,
  0.0004299959, -0.0016043, -0.004559465, -0.0009546667, -4.66862e-05, 
    4.66862e-05, 0.0009546667, 0.004559465, 0.0016043, -0.0004299959,
  0.0004299959, -0.0016043, -0.004559465, -0.0009546667, -4.66862e-05, 
    4.66862e-05, 0.0009546667, 0.004559465, 0.0016043, -0.0004299959,
  0.0002650476, -0.0009887358, -0.004477448, -0.002047871, -0.0003399205, 
    0.0003399205, 0.002047871, 0.004477448, 0.0009887358, -0.0002650476,
  0, -0.0001630833, -0.004002416, -0.002663461, -0.0008098975, 0.0008098975, 
    0.002663461, 0.004002416, 0.0001630833, 0,
  0, 0, 2.959485e-06, -4.599014e-05, -4.764587e-05, 4.764587e-05, 
    4.599014e-05, -2.959485e-06, 0, 0,
  0, 0, 0, 1.179233e-05, 1.274914e-05, -1.274914e-05, -1.179233e-05, 0, 0, 0,
  0, 0, 0, 7.582334e-06, 8.342955e-06, -8.342955e-06, -7.582334e-06, 0, 0, 0,
  0, 0, 9.544734e-06, -2.920879e-05, -3.116686e-05, 3.116686e-05, 
    2.920879e-05, -9.544734e-06, 0, 0,
  0, -9.885567e-05, -0.002666362, -0.001774951, -0.0005401318, 0.0005401318, 
    0.001774951, 0.002666362, 9.885567e-05, 0,
  0.0001743191, -0.0006503563, -0.00298789, -0.001356395, -0.0002240145, 
    0.0002240145, 0.001356395, 0.00298789, 0.0006503563, -0.0001743191,
  0.0002834205, -0.001057508, -0.003044778, -0.0006273668, -3.050758e-05, 
    3.050758e-05, 0.0006273668, 0.003044778, 0.001057508, -0.0002834205,
  0.0002834205, -0.001057508, -0.003044778, -0.0006273668, -3.050758e-05, 
    3.050758e-05, 0.0006273668, 0.003044778, 0.001057508, -0.0002834205,
  0.0001743191, -0.0006503563, -0.00298789, -0.001356395, -0.0002240145, 
    0.0002240145, 0.001356395, 0.00298789, 0.0006503563, -0.0001743191,
  0, -9.885567e-05, -0.002666362, -0.001774951, -0.0005401318, 0.0005401318, 
    0.001774951, 0.002666362, 9.885567e-05, 0,
  0, 0, 9.544734e-06, -2.920879e-05, -3.116686e-05, 3.116686e-05, 
    2.920879e-05, -9.544734e-06, 0, 0,
  0, 0, 0, 7.582334e-06, 8.342955e-06, -8.342955e-06, -7.582334e-06, 0, 0, 0,
  0, 0, 0, 3.613859e-06, 4.069061e-06, -4.069061e-06, -3.613859e-06, 0, 0, 0,
  0, 0, 8.185861e-06, -1.373546e-05, -1.519242e-05, 1.519242e-05, 
    1.373546e-05, -8.185861e-06, 0, 0,
  0, -4.47583e-05, -0.001324375, -0.000883024, -0.0002690957, 0.0002690957, 
    0.000883024, 0.001324375, 4.47583e-05, 0,
  8.544845e-05, -0.0003188381, -0.001488222, -0.0006720317, -0.0001104672, 
    0.0001104672, 0.0006720317, 0.001488222, 0.0003188381, -8.544845e-05,
  0.0001391938, -0.0005194148, -0.001518787, -0.0003086543, -1.501882e-05, 
    1.501882e-05, 0.0003086543, 0.001518787, 0.0005194148, -0.0001391938,
  0.0001391938, -0.0005194148, -0.001518787, -0.0003086543, -1.501882e-05, 
    1.501882e-05, 0.0003086543, 0.001518787, 0.0005194148, -0.0001391938,
  8.544845e-05, -0.0003188381, -0.001488222, -0.0006720317, -0.0001104672, 
    0.0001104672, 0.0006720317, 0.001488222, 0.0003188381, -8.544845e-05,
  0, -4.47583e-05, -0.001324375, -0.000883024, -0.0002690957, 0.0002690957, 
    0.000883024, 0.001324375, 4.47583e-05, 0,
  0, 0, 8.185861e-06, -1.373546e-05, -1.519242e-05, 1.519242e-05, 
    1.373546e-05, -8.185861e-06, 0, 0,
  0, 0, 0, 3.613859e-06, 4.069061e-06, -4.069061e-06, -3.613859e-06, 0, 0, 0,
  0, 0, 0, 5.861484e-10, 3.122964e-10, -3.122964e-10, -5.861484e-10, 0, 0, 0,
  0, 0, -1.156787e-08, -4.258139e-09, -1.098778e-09, 1.098778e-09, 
    4.258139e-09, 1.156787e-08, 0, 0,
  0, -1.331484e-08, -2.344673e-08, -1.553574e-08, -4.864146e-09, 
    4.864146e-09, 1.553574e-08, 2.344673e-08, 1.331484e-08, 0,
  5.822006e-09, -2.387134e-08, -2.44924e-08, -1.537197e-08, -5.10307e-09, 
    5.10307e-09, 1.537197e-08, 2.44924e-08, 2.387134e-08, -5.822006e-09,
  7.003699e-09, -2.873023e-08, -2.523416e-08, -1.533583e-08, -5.883404e-09, 
    5.883404e-09, 1.533583e-08, 2.523416e-08, 2.873023e-08, -7.003699e-09,
  7.003699e-09, -2.873023e-08, -2.523416e-08, -1.533583e-08, -5.883404e-09, 
    5.883404e-09, 1.533583e-08, 2.523416e-08, 2.873023e-08, -7.003699e-09,
  5.822006e-09, -2.387134e-08, -2.44924e-08, -1.537197e-08, -5.10307e-09, 
    5.10307e-09, 1.537197e-08, 2.44924e-08, 2.387134e-08, -5.822006e-09,
  0, -1.331484e-08, -2.344673e-08, -1.553574e-08, -4.864146e-09, 
    4.864146e-09, 1.553574e-08, 2.344673e-08, 1.331484e-08, 0,
  0, 0, -1.156787e-08, -4.258139e-09, -1.098778e-09, 1.098778e-09, 
    4.258139e-09, 1.156787e-08, 0, 0,
  0, 0, 0, 5.861484e-10, 3.122964e-10, -3.122964e-10, -5.861484e-10, 0, 0, 0,
  0, 0, 0, 3.446963e-05, 2.833646e-05, -2.833646e-05, -3.446963e-05, 0, 0, 0,
  0, 0, -0.0002989912, -0.0001408909, -0.0001062195, 0.0001062195, 
    0.0001408909, 0.0002989912, 0, 0,
  0, -0.000761056, -0.008313667, -0.005538933, -0.001694023, 0.001694023, 
    0.005538933, 0.008313667, 0.000761056, 0,
  0.0006145203, -0.002291939, -0.009221511, -0.004532514, -0.0008527749, 
    0.0008527749, 0.004532514, 0.009221511, 0.002291939, -0.0006145203,
  0.0009423745, -0.003524209, -0.009451356, -0.002400297, -0.0001504265, 
    0.0001504265, 0.002400297, 0.009451356, 0.003524209, -0.0009423745,
  0.0009423745, -0.003524209, -0.009451356, -0.002400297, -0.0001504265, 
    0.0001504265, 0.002400297, 0.009451356, 0.003524209, -0.0009423745,
  0.0006145203, -0.002291939, -0.009221511, -0.004532514, -0.0008527749, 
    0.0008527749, 0.004532514, 0.009221511, 0.002291939, -0.0006145203,
  0, -0.000761056, -0.008313667, -0.005538933, -0.001694023, 0.001694023, 
    0.005538933, 0.008313667, 0.000761056, 0,
  0, 0, -0.0002989912, -0.0001408909, -0.0001062195, 0.0001062195, 
    0.0001408909, 0.0002989912, 0, 0,
  0, 0, 0, 3.446963e-05, 2.833646e-05, -2.833646e-05, -3.446963e-05, 0, 0, 0,
  0, 0, 0, 3.265457e-05, 2.809974e-05, -2.809974e-05, -3.265457e-05, 0, 0, 0,
  0, 0, -0.0002554863, -0.0001338267, -0.0001052244, 0.0001052244, 
    0.0001338267, 0.0002554863, 0, 0,
  0, -0.0006946157, -0.008243145, -0.005477678, -0.001671177, 0.001671177, 
    0.005477678, 0.008243145, 0.0006946157, 0,
  0.0006018683, -0.002244339, -0.009120974, -0.004456076, -0.0008233186, 
    0.0008233186, 0.004456076, 0.009120974, 0.002244339, -0.0006018683,
  0.0009309254, -0.003476808, -0.009326496, -0.002324953, -0.0001416827, 
    0.0001416827, 0.002324953, 0.009326496, 0.003476808, -0.0009309254,
  0.0009309254, -0.003476808, -0.009326496, -0.002324953, -0.0001416827, 
    0.0001416827, 0.002324953, 0.009326496, 0.003476808, -0.0009309254,
  0.0006018683, -0.002244339, -0.009120974, -0.004456076, -0.0008233186, 
    0.0008233186, 0.004456076, 0.009120974, 0.002244339, -0.0006018683,
  0, -0.0006946157, -0.008243145, -0.005477678, -0.001671177, 0.001671177, 
    0.005477678, 0.008243145, 0.0006946157, 0,
  0, 0, -0.0002554863, -0.0001338267, -0.0001052244, 0.0001052244, 
    0.0001338267, 0.0002554863, 0, 0,
  0, 0, 0, 3.265457e-05, 2.809974e-05, -2.809974e-05, -3.265457e-05, 0, 0, 0,
  0, 0, 0, 2.965407e-05, 2.726686e-05, -2.726686e-05, -2.965407e-05, 0, 0, 0,
  0, 0, -0.0001762706, -0.0001208219, -0.0001019677, 0.0001019677, 
    0.0001208219, 0.0001762706, 0, 0,
  0, -0.0005744161, -0.007975801, -0.005282386, -0.001603614, 0.001603614, 
    0.005282386, 0.007975801, 0.0005744161, 0,
  0.000569397, -0.002123483, -0.008808539, -0.004224174, -0.0007551908, 
    0.0007551908, 0.004224174, 0.008808539, 0.002123483, -0.000569397,
  0.0008949178, -0.003339963, -0.008962623, -0.002135323, -0.0001242063, 
    0.0001242063, 0.002135323, 0.008962623, 0.003339963, -0.0008949178,
  0.0008949178, -0.003339963, -0.008962623, -0.002135323, -0.0001242063, 
    0.0001242063, 0.002135323, 0.008962623, 0.003339963, -0.0008949178,
  0.000569397, -0.002123483, -0.008808539, -0.004224174, -0.0007551908, 
    0.0007551908, 0.004224174, 0.008808539, 0.002123483, -0.000569397,
  0, -0.0005744161, -0.007975801, -0.005282386, -0.001603614, 0.001603614, 
    0.005282386, 0.007975801, 0.0005744161, 0,
  0, 0, -0.0001762706, -0.0001208219, -0.0001019677, 0.0001019677, 
    0.0001208219, 0.0001762706, 0, 0,
  0, 0, 0, 2.965407e-05, 2.726686e-05, -2.726686e-05, -2.965407e-05, 0, 0, 0,
  0, 0, 0, 2.58518e-05, 2.493356e-05, -2.493356e-05, -2.58518e-05, 0, 0, 0,
  0, 0, -0.0001073958, -0.0001042298, -9.322522e-05, 9.322522e-05, 
    0.0001042298, 0.0001073958, 0, 0,
  0, -0.0004545368, -0.007372889, -0.00488117, -0.001478728, 0.001478728, 
    0.00488117, 0.007372889, 0.0004545368, 0,
  0.0005155338, -0.001922653, -0.008155355, -0.003846478, -0.0006677705, 
    0.0006677705, 0.003846478, 0.008155355, 0.001922653, -0.0005155338,
  0.0008197739, -0.003058663, -0.008276966, -0.001887635, -0.000103518, 
    0.000103518, 0.001887635, 0.008276966, 0.003058663, -0.0008197739,
  0.0008197739, -0.003058663, -0.008276966, -0.001887635, -0.000103518, 
    0.000103518, 0.001887635, 0.008276966, 0.003058663, -0.0008197739,
  0.0005155338, -0.001922653, -0.008155355, -0.003846478, -0.0006677705, 
    0.0006677705, 0.003846478, 0.008155355, 0.001922653, -0.0005155338,
  0, -0.0004545368, -0.007372889, -0.00488117, -0.001478728, 0.001478728, 
    0.00488117, 0.007372889, 0.0004545368, 0,
  0, 0, -0.0001073958, -0.0001042298, -9.322522e-05, 9.322522e-05, 
    0.0001042298, 0.0001073958, 0, 0,
  0, 0, 0, 2.58518e-05, 2.493356e-05, -2.493356e-05, -2.58518e-05, 0, 0, 0,
  0, 0, 0, 2.146614e-05, 2.142994e-05, -2.142994e-05, -2.146614e-05, 0, 0, 0,
  0, 0, -5.649689e-05, -8.555062e-05, -8.012012e-05, 8.012012e-05, 
    8.555062e-05, 5.649689e-05, 0, 0,
  0, -0.0003462129, -0.006446572, -0.004270537, -0.00129395, 0.00129395, 
    0.004270537, 0.006446572, 0.0003462129, 0,
  0.0004427115, -0.001651167, -0.007149083, -0.003329981, -0.0005673318, 
    0.0005673318, 0.003329981, 0.007149083, 0.001651167, -0.0004427115,
  0.0007094275, -0.002646727, -0.007253477, -0.001600625, -8.340323e-05, 
    8.340323e-05, 0.001600625, 0.007253477, 0.002646727, -0.0007094275,
  0.0007094275, -0.002646727, -0.007253477, -0.001600625, -8.340323e-05, 
    8.340323e-05, 0.001600625, 0.007253477, 0.002646727, -0.0007094275,
  0.0004427115, -0.001651167, -0.007149083, -0.003329981, -0.0005673318, 
    0.0005673318, 0.003329981, 0.007149083, 0.001651167, -0.0004427115,
  0, -0.0003462129, -0.006446572, -0.004270537, -0.00129395, 0.00129395, 
    0.004270537, 0.006446572, 0.0003462129, 0,
  0, 0, -5.649689e-05, -8.555062e-05, -8.012012e-05, 8.012012e-05, 
    8.555062e-05, 5.649689e-05, 0, 0,
  0, 0, 0, 2.146614e-05, 2.142994e-05, -2.142994e-05, -2.146614e-05, 0, 0, 0,
  0, 0, 0, 1.685587e-05, 1.727621e-05, -1.727621e-05, -1.685587e-05, 0, 0, 0,
  0, 0, -2.242266e-05, -6.639662e-05, -6.457946e-05, 6.457946e-05, 
    6.639662e-05, 2.242266e-05, 0, 0,
  0, -0.0002518299, -0.005292843, -0.003508329, -0.001063868, 0.001063868, 
    0.003508329, 0.005292843, 0.0002518299, 0,
  0.0003578071, -0.001334621, -0.005883555, -0.002713289, -0.0004570856, 
    0.0004570856, 0.002713289, 0.005883555, 0.001334621, -0.0003578071,
  0.0005763965, -0.002150422, -0.005972451, -0.001286073, -6.48932e-05, 
    6.48932e-05, 0.001286073, 0.005972451, 0.002150422, -0.0005763965,
  0.0005763965, -0.002150422, -0.005972451, -0.001286073, -6.48932e-05, 
    6.48932e-05, 0.001286073, 0.005972451, 0.002150422, -0.0005763965,
  0.0003578071, -0.001334621, -0.005883555, -0.002713289, -0.0004570856, 
    0.0004570856, 0.002713289, 0.005883555, 0.001334621, -0.0003578071,
  0, -0.0002518299, -0.005292843, -0.003508329, -0.001063868, 0.001063868, 
    0.003508329, 0.005292843, 0.0002518299, 0,
  0, 0, -2.242266e-05, -6.639662e-05, -6.457946e-05, 6.457946e-05, 
    6.639662e-05, 2.242266e-05, 0, 0,
  0, 0, 0, 1.685587e-05, 1.727621e-05, -1.727621e-05, -1.685587e-05, 0, 0, 0,
  0, 0, 0, 1.229173e-05, 1.285302e-05, -1.285302e-05, -1.229173e-05, 0, 0, 0,
  0, 0, -2.790395e-06, -4.78558e-05, -4.803204e-05, 4.803204e-05, 
    4.78558e-05, 2.790395e-06, 0, 0,
  0, -0.0001719668, -0.004010062, -0.002658849, -0.0008069191, 0.0008069191, 
    0.002658849, 0.004010062, 0.0001719668, 0,
  0.0002673276, -0.0009972363, -0.004465958, -0.002041946, -0.0003415819, 
    0.0003415819, 0.002041946, 0.004465958, 0.0009972363, -0.0002673276,
  0.0004321113, -0.001612196, -0.004536331, -0.0009582682, -4.758104e-05, 
    4.758104e-05, 0.0009582682, 0.004536331, 0.001612196, -0.0004321113,
  0.0004321113, -0.001612196, -0.004536331, -0.0009582682, -4.758104e-05, 
    4.758104e-05, 0.0009582682, 0.004536331, 0.001612196, -0.0004321113,
  0.0002673276, -0.0009972363, -0.004465958, -0.002041946, -0.0003415819, 
    0.0003415819, 0.002041946, 0.004465958, 0.0009972363, -0.0002673276,
  0, -0.0001719668, -0.004010062, -0.002658849, -0.0008069191, 0.0008069191, 
    0.002658849, 0.004010062, 0.0001719668, 0,
  0, 0, -2.790395e-06, -4.78558e-05, -4.803204e-05, 4.803204e-05, 
    4.78558e-05, 2.790395e-06, 0, 0,
  0, 0, 0, 1.229173e-05, 1.285302e-05, -1.285302e-05, -1.229173e-05, 0, 0, 0,
  0, 0, 0, 7.908131e-06, 8.413174e-06, -8.413174e-06, -7.908131e-06, 0, 0, 0,
  0, 0, 5.767954e-06, -3.042558e-05, -3.142826e-05, 3.142826e-05, 
    3.042558e-05, -5.767954e-06, 0, 0,
  0, -0.0001047961, -0.002672944, -0.001772953, -0.000538476, 0.000538476, 
    0.001772953, 0.002672944, 0.0001047961, 0,
  0.0001758832, -0.0006561888, -0.002982057, -0.00135321, -0.0002252401, 
    0.0002252401, 0.00135321, 0.002982057, 0.0006561888, -0.0001758832,
  0.0002848972, -0.001063018, -0.003031253, -0.0006300837, -3.111303e-05, 
    3.111303e-05, 0.0006300837, 0.003031253, 0.001063018, -0.0002848972,
  0.0002848972, -0.001063018, -0.003031253, -0.0006300837, -3.111303e-05, 
    3.111303e-05, 0.0006300837, 0.003031253, 0.001063018, -0.0002848972,
  0.0001758832, -0.0006561888, -0.002982057, -0.00135321, -0.0002252401, 
    0.0002252401, 0.00135321, 0.002982057, 0.0006561888, -0.0001758832,
  0, -0.0001047961, -0.002672944, -0.001772953, -0.000538476, 0.000538476, 
    0.001772953, 0.002672944, 0.0001047961, 0,
  0, 0, 5.767954e-06, -3.042558e-05, -3.142826e-05, 3.142826e-05, 
    3.042558e-05, -5.767954e-06, 0, 0,
  0, 0, 0, 7.908131e-06, 8.413174e-06, -8.413174e-06, -7.908131e-06, 0, 0, 0,
  0, 0, 0, 3.767081e-06, 4.104208e-06, -4.104208e-06, -3.767081e-06, 0, 0, 0,
  0, 0, 6.41051e-06, -1.430753e-05, -1.532345e-05, 1.532345e-05, 
    1.430753e-05, -6.41051e-06, 0, 0,
  0, -4.760958e-05, -0.001328308, -0.0008826931, -0.000268516, 0.000268516, 
    0.0008826931, 0.001328308, 4.760958e-05, 0,
  8.623255e-05, -0.000321763, -0.001486439, -0.0006711513, -0.0001111782, 
    0.0001111782, 0.0006711513, 0.001486439, 0.000321763, -8.623255e-05,
  0.0001399608, -0.0005222771, -0.001513435, -0.0003103066, -1.533146e-05, 
    1.533146e-05, 0.0003103066, 0.001513435, 0.0005222771, -0.0001399608,
  0.0001399608, -0.0005222771, -0.001513435, -0.0003103066, -1.533146e-05, 
    1.533146e-05, 0.0003103066, 0.001513435, 0.0005222771, -0.0001399608,
  8.623255e-05, -0.000321763, -0.001486439, -0.0006711513, -0.0001111782, 
    0.0001111782, 0.0006711513, 0.001486439, 0.000321763, -8.623255e-05,
  0, -4.760958e-05, -0.001328308, -0.0008826931, -0.000268516, 0.000268516, 
    0.0008826931, 0.001328308, 4.760958e-05, 0,
  0, 0, 6.41051e-06, -1.430753e-05, -1.532345e-05, 1.532345e-05, 
    1.430753e-05, -6.41051e-06, 0, 0,
  0, 0, 0, 3.767081e-06, 4.104208e-06, -4.104208e-06, -3.767081e-06, 0, 0, 0,
  0, 0, 0, 5.863201e-10, 3.123937e-10, -3.123937e-10, -5.863201e-10, 0, 0, 0,
  0, 0, -1.158092e-08, -4.263859e-09, -1.099315e-09, 1.099315e-09, 
    4.263859e-09, 1.158092e-08, 0, 0,
  0, -1.334284e-08, -2.343999e-08, -1.552301e-08, -4.861426e-09, 
    4.861426e-09, 1.552301e-08, 2.343999e-08, 1.334284e-08, 0,
  5.82523e-09, -2.390036e-08, -2.44425e-08, -1.535468e-08, -5.105515e-09, 
    5.105515e-09, 1.535468e-08, 2.44425e-08, 2.390036e-08, -5.82523e-09,
  7.004086e-09, -2.875323e-08, -2.516461e-08, -1.534258e-08, -5.903839e-09, 
    5.903839e-09, 1.534258e-08, 2.516461e-08, 2.875323e-08, -7.004086e-09,
  7.004086e-09, -2.875323e-08, -2.516461e-08, -1.534258e-08, -5.903839e-09, 
    5.903839e-09, 1.534258e-08, 2.516461e-08, 2.875323e-08, -7.004086e-09,
  5.82523e-09, -2.390036e-08, -2.44425e-08, -1.535468e-08, -5.105515e-09, 
    5.105515e-09, 1.535468e-08, 2.44425e-08, 2.390036e-08, -5.82523e-09,
  0, -1.334284e-08, -2.343999e-08, -1.552301e-08, -4.861426e-09, 
    4.861426e-09, 1.552301e-08, 2.343999e-08, 1.334284e-08, 0,
  0, 0, -1.158092e-08, -4.263859e-09, -1.099315e-09, 1.099315e-09, 
    4.263859e-09, 1.158092e-08, 0, 0,
  0, 0, 0, 5.863201e-10, 3.123937e-10, -3.123937e-10, -5.863201e-10, 0, 0, 0,
  0, 0, 0, 4.86494e-05, 2.325717e-05, -2.325717e-05, -4.86494e-05, 0, 0, 0,
  0, -0.000122941, 0.0005033952, -0.0001888947, -8.905558e-05, 8.905558e-05, 
    0.0001888947, -0.0005033952, 0.000122941, 0,
  0, 0.0005770404, -0.002340529, -0.005456394, -0.001691033, 0.001691033, 
    0.005456394, 0.002340529, -0.0005770404, 0,
  0.0005071253, -0.001891851, -0.008948468, -0.004253624, -0.0008928971, 
    0.0008928971, 0.004253624, 0.008948468, 0.001891851, -0.0005071253,
  0.0009713179, -0.003632271, -0.00943802, -0.002438161, -0.0001476524, 
    0.0001476524, 0.002438161, 0.00943802, 0.003632271, -0.0009713179,
  0.0009713179, -0.003632271, -0.00943802, -0.002438161, -0.0001476524, 
    0.0001476524, 0.002438161, 0.00943802, 0.003632271, -0.0009713179,
  0.0005071253, -0.001891851, -0.008948468, -0.004253624, -0.0008928971, 
    0.0008928971, 0.004253624, 0.008948468, 0.001891851, -0.0005071253,
  0, 0.0005770404, -0.002340529, -0.005456394, -0.001691033, 0.001691033, 
    0.005456394, 0.002340529, -0.0005770404, 0,
  0, -0.000122941, 0.0005033952, -0.0001888947, -8.905558e-05, 8.905558e-05, 
    0.0001888947, -0.0005033952, 0.000122941, 0,
  0, 0, 0, 4.86494e-05, 2.325717e-05, -2.325717e-05, -4.86494e-05, 0, 0, 0,
  0, 0, 0, 4.504287e-05, 2.358981e-05, -2.358981e-05, -4.504287e-05, 0, 0, 0,
  0, -0.0001251832, 0.0005016397, -0.0001763244, -8.975093e-05, 8.975093e-05, 
    0.0001763244, -0.0005016397, 0.0001251832, 0,
  0, 0.0005752536, -0.002295947, -0.005395042, -0.001668034, 0.001668034, 
    0.005395042, 0.002295947, -0.0005752536, 0,
  0.000493344, -0.001841575, -0.008847, -0.004195032, -0.0008596442, 
    0.0008596442, 0.004195032, 0.008847, 0.001841575, -0.000493344,
  0.0009601261, -0.003585364, -0.00931478, -0.002360326, -0.0001393442, 
    0.0001393442, 0.002360326, 0.00931478, 0.003585364, -0.0009601261,
  0.0009601261, -0.003585364, -0.00931478, -0.002360326, -0.0001393442, 
    0.0001393442, 0.002360326, 0.00931478, 0.003585364, -0.0009601261,
  0.000493344, -0.001841575, -0.008847, -0.004195032, -0.0008596442, 
    0.0008596442, 0.004195032, 0.008847, 0.001841575, -0.000493344,
  0, 0.0005752536, -0.002295947, -0.005395042, -0.001668034, 0.001668034, 
    0.005395042, 0.002295947, -0.0005752536, 0,
  0, -0.0001251832, 0.0005016397, -0.0001763244, -8.975093e-05, 8.975093e-05, 
    0.0001763244, -0.0005016397, 0.0001251832, 0,
  0, 0, 0, 4.504287e-05, 2.358981e-05, -2.358981e-05, -4.504287e-05, 0, 0, 0,
  0, 0, 0, 3.923894e-05, 2.362618e-05, -2.362618e-05, -3.923894e-05, 0, 0, 0,
  0, -0.0001248465, 0.0004885047, -0.0001540941, -8.927784e-05, 8.927784e-05, 
    0.0001540941, -0.0004885047, 0.0001248465, 0,
  0, 0.0005574753, -0.002183635, -0.005204882, -0.001599355, 0.001599355, 
    0.005204882, 0.002183635, -0.0005574753, 0,
  0.0004607817, -0.001720755, -0.00853559, -0.003996574, -0.0007861073, 
    0.0007861073, 0.003996574, 0.00853559, 0.001720755, -0.0004607817,
  0.000924008, -0.003447955, -0.008954303, -0.00216685, -0.0001223268, 
    0.0001223268, 0.00216685, 0.008954303, 0.003447955, -0.000924008,
  0.000924008, -0.003447955, -0.008954303, -0.00216685, -0.0001223268, 
    0.0001223268, 0.00216685, 0.008954303, 0.003447955, -0.000924008,
  0.0004607817, -0.001720755, -0.00853559, -0.003996574, -0.0007861073, 
    0.0007861073, 0.003996574, 0.00853559, 0.001720755, -0.0004607817,
  0, 0.0005574753, -0.002183635, -0.005204882, -0.001599355, 0.001599355, 
    0.005204882, 0.002183635, -0.0005574753, 0,
  0, -0.0001248465, 0.0004885047, -0.0001540941, -8.927784e-05, 8.927784e-05, 
    0.0001540941, -0.0004885047, 0.0001248465, 0,
  0, 0, 0, 3.923894e-05, 2.362618e-05, -2.362618e-05, -3.923894e-05, 0, 0, 0,
  0, 0, 0, 3.298846e-05, 2.209667e-05, -2.209667e-05, -3.298846e-05, 0, 0, 0,
  0, -0.0001174738, 0.0004535116, -0.0001292149, -8.322528e-05, 8.322528e-05, 
    0.0001292149, -0.0004535116, 0.0001174738, 0,
  0, 0.000513422, -0.001988313, -0.004817074, -0.001472444, 0.001472444, 
    0.004817074, 0.001988313, -0.000513422, 0,
  0.0004127499, -0.001541335, -0.007900783, -0.003653675, -0.0006939937, 
    0.0006939937, 0.003653675, 0.007900783, 0.001541335, -0.0004127499,
  0.0008472838, -0.003160817, -0.00827109, -0.001915359, -0.0001019367, 
    0.0001019367, 0.001915359, 0.00827109, 0.003160817, -0.0008472838,
  0.0008472838, -0.003160817, -0.00827109, -0.001915359, -0.0001019367, 
    0.0001019367, 0.001915359, 0.00827109, 0.003160817, -0.0008472838,
  0.0004127499, -0.001541335, -0.007900783, -0.003653675, -0.0006939937, 
    0.0006939937, 0.003653675, 0.007900783, 0.001541335, -0.0004127499,
  0, 0.000513422, -0.001988313, -0.004817074, -0.001472444, 0.001472444, 
    0.004817074, 0.001988313, -0.000513422, 0,
  0, -0.0001174738, 0.0004535116, -0.0001292149, -8.322528e-05, 8.322528e-05, 
    0.0001292149, -0.0004535116, 0.0001174738, 0,
  0, 0, 0, 3.298846e-05, 2.209667e-05, -2.209667e-05, -3.298846e-05, 0, 0, 0,
  0, 0, 0, 2.664342e-05, 1.928389e-05, -1.928389e-05, -2.664342e-05, 0, 0, 0,
  0, -0.0001035608, 0.0003970476, -0.0001038137, -7.248516e-05, 7.248516e-05, 
    0.0001038137, -0.0003970476, 0.0001035608, 0,
  0, 0.0004460113, -0.001716495, -0.004223715, -0.001285968, 0.001285968, 
    0.004223715, 0.001716495, -0.0004460113, 0,
  0.000351859, -0.001313798, -0.006928134, -0.003172668, -0.0005888975, 
    0.0005888975, 0.003172668, 0.006928134, 0.001313798, -0.000351859,
  0.0007338061, -0.002737319, -0.007249506, -0.00162399, -8.213058e-05, 
    8.213058e-05, 0.00162399, 0.007249506, 0.002737319, -0.0007338061,
  0.0007338061, -0.002737319, -0.007249506, -0.00162399, -8.213058e-05, 
    8.213058e-05, 0.00162399, 0.007249506, 0.002737319, -0.0007338061,
  0.000351859, -0.001313798, -0.006928134, -0.003172668, -0.0005888975, 
    0.0005888975, 0.003172668, 0.006928134, 0.001313798, -0.000351859,
  0, 0.0004460113, -0.001716495, -0.004223715, -0.001285968, 0.001285968, 
    0.004223715, 0.001716495, -0.0004460113, 0,
  0, -0.0001035608, 0.0003970476, -0.0001038137, -7.248516e-05, 7.248516e-05, 
    0.0001038137, -0.0003970476, 0.0001035608, 0,
  0, 0, 0, 2.664342e-05, 1.928389e-05, -1.928389e-05, -2.664342e-05, 0, 0, 0,
  0, 0, 0, 2.044338e-05, 1.572823e-05, -1.572823e-05, -2.044338e-05, 0, 0, 0,
  0, -8.528172e-05, 0.0003256902, -7.914679e-05, -5.902622e-05, 5.902622e-05, 
    7.914679e-05, -0.0003256902, 8.528172e-05, 0,
  0, 0.0003635667, -0.001394031, -0.00347805, -0.001055357, 0.001055357, 
    0.00347805, 0.001394031, -0.0003635667, 0,
  0.0002829162, -0.001056253, -0.005705225, -0.002591366, -0.000473982, 
    0.000473982, 0.002591366, 0.005705225, 0.001056253, -0.0002829162,
  0.0005965838, -0.0022255, -0.005970362, -0.001304716, -6.393938e-05, 
    6.393938e-05, 0.001304716, 0.005970362, 0.0022255, -0.0005965838,
  0.0005965838, -0.0022255, -0.005970362, -0.001304716, -6.393938e-05, 
    6.393938e-05, 0.001304716, 0.005970362, 0.0022255, -0.0005965838,
  0.0002829162, -0.001056253, -0.005705225, -0.002591366, -0.000473982, 
    0.000473982, 0.002591366, 0.005705225, 0.001056253, -0.0002829162,
  0, 0.0003635667, -0.001394031, -0.00347805, -0.001055357, 0.001055357, 
    0.00347805, 0.001394031, -0.0003635667, 0,
  0, -8.528172e-05, 0.0003256902, -7.914679e-05, -5.902622e-05, 5.902622e-05, 
    7.914679e-05, -0.0003256902, 8.528172e-05, 0,
  0, 0, 0, 2.044338e-05, 1.572823e-05, -1.572823e-05, -2.044338e-05, 0, 0, 0,
  0, 0, 0, 1.460284e-05, 1.181465e-05, -1.181465e-05, -1.460284e-05, 0, 0, 0,
  0, -6.459056e-05, 0.0002460892, -5.613481e-05, -4.427704e-05, 4.427704e-05, 
    5.613481e-05, -0.0002460892, 6.459056e-05, 0,
  0, 0.0002734499, -0.001046096, -0.002642252, -0.0007992044, 0.0007992044, 
    0.002642252, 0.001046096, -0.0002734499, 0,
  0.0002105939, -0.0007861596, -0.004334302, -0.001954187, -0.0003539496, 
    0.0003539496, 0.001954187, 0.004334302, 0.0007861596, -0.0002105939,
  0.000447504, -0.001669488, -0.004536202, -0.0009721543, -4.692788e-05, 
    4.692788e-05, 0.0009721543, 0.004536202, 0.001669488, -0.000447504,
  0.000447504, -0.001669488, -0.004536202, -0.0009721543, -4.692788e-05, 
    4.692788e-05, 0.0009721543, 0.004536202, 0.001669488, -0.000447504,
  0.0002105939, -0.0007861596, -0.004334302, -0.001954187, -0.0003539496, 
    0.0003539496, 0.001954187, 0.004334302, 0.0007861596, -0.0002105939,
  0, 0.0002734499, -0.001046096, -0.002642252, -0.0007992044, 0.0007992044, 
    0.002642252, 0.001046096, -0.0002734499, 0,
  0, -6.459056e-05, 0.0002460892, -5.613481e-05, -4.427704e-05, 4.427704e-05, 
    5.613481e-05, -0.0002460892, 6.459056e-05, 0,
  0, 0, 0, 1.460284e-05, 1.181465e-05, -1.181465e-05, -1.460284e-05, 0, 0, 0,
  0, 0, 0, 9.211845e-06, 7.80042e-06, -7.80042e-06, -9.211845e-06, 0, 0, 0,
  0, -4.292298e-05, 0.0001632886, -3.513769e-05, -2.919402e-05, 2.919402e-05, 
    3.513769e-05, -0.0001632886, 4.292298e-05, 0,
  0, 0.0001808726, -0.0006909294, -0.00176618, -0.0005327126, 0.0005327126, 
    0.00176618, 0.0006909294, -0.0001808726, 0,
  0.0001381627, -0.0005157209, -0.00289724, -0.001297592, -0.0002333162, 
    0.0002333162, 0.001297592, 0.00289724, 0.0005157209, -0.0001381627,
  0.0002952171, -0.00110146, -0.003032865, -0.0006393747, -3.072609e-05, 
    3.072609e-05, 0.0006393747, 0.003032865, 0.00110146, -0.0002952171,
  0.0002952171, -0.00110146, -0.003032865, -0.0006393747, -3.072609e-05, 
    3.072609e-05, 0.0006393747, 0.003032865, 0.00110146, -0.0002952171,
  0.0001381627, -0.0005157209, -0.00289724, -0.001297592, -0.0002333162, 
    0.0002333162, 0.001297592, 0.00289724, 0.0005157209, -0.0001381627,
  0, 0.0001808726, -0.0006909294, -0.00176618, -0.0005327126, 0.0005327126, 
    0.00176618, 0.0006909294, -0.0001808726, 0,
  0, -4.292298e-05, 0.0001632886, -3.513769e-05, -2.919402e-05, 2.919402e-05, 
    3.513769e-05, -0.0001632886, 4.292298e-05, 0,
  0, 0, 0, 9.211845e-06, 7.80042e-06, -7.80042e-06, -9.211845e-06, 0, 0, 0,
  0, 0, 0, 4.301308e-06, 3.837732e-06, -3.837732e-06, -4.301308e-06, 0, 0, 0,
  0, -2.121002e-05, 8.059232e-05, -1.626051e-05, -1.434243e-05, 1.434243e-05, 
    1.626051e-05, -8.059232e-05, 2.121002e-05, 0,
  0, 8.90798e-05, -0.0003399263, -0.0008812804, -0.0002654715, 0.0002654715, 
    0.0008812804, 0.0003399263, -8.90798e-05, 0,
  6.754683e-05, -0.0002521111, -0.00144566, -0.0006449149, -0.0001151896, 
    0.0001151896, 0.0006449149, 0.00144566, 0.0002521111, -6.754683e-05,
  0.0001451101, -0.0005414747, -0.001515442, -0.0003151101, -1.516404e-05, 
    1.516404e-05, 0.0003151101, 0.001515442, 0.0005414747, -0.0001451101,
  0.0001451101, -0.0005414747, -0.001515442, -0.0003151101, -1.516404e-05, 
    1.516404e-05, 0.0003151101, 0.001515442, 0.0005414747, -0.0001451101,
  6.754683e-05, -0.0002521111, -0.00144566, -0.0006449149, -0.0001151896, 
    0.0001151896, 0.0006449149, 0.00144566, 0.0002521111, -6.754683e-05,
  0, 8.90798e-05, -0.0003399263, -0.0008812804, -0.0002654715, 0.0002654715, 
    0.0008812804, 0.0003399263, -8.90798e-05, 0,
  0, -2.121002e-05, 8.059232e-05, -1.626051e-05, -1.434243e-05, 1.434243e-05, 
    1.626051e-05, -8.059232e-05, 2.121002e-05, 0,
  0, 0, 0, 4.301308e-06, 3.837732e-06, -3.837732e-06, -4.301308e-06, 0, 0, 0,
  0, 0, 0, 8.882792e-10, 2.049165e-10, -2.049165e-10, -8.882792e-10, 0, 0, 0,
  0, 2.319781e-09, -4.599584e-09, -4.862396e-09, -9.173195e-10, 9.173195e-10, 
    4.862396e-09, 4.599584e-09, -2.319781e-09, 0,
  0, -4.230289e-09, -1.879162e-08, -1.511646e-08, -4.975775e-09, 
    4.975775e-09, 1.511646e-08, 1.879162e-08, 4.230289e-09, 0,
  5.804671e-09, -2.381888e-08, -2.450905e-08, -1.50993e-08, -5.1423e-09, 
    5.1423e-09, 1.50993e-08, 2.450905e-08, 2.381888e-08, -5.804671e-09,
  7.008032e-09, -2.878978e-08, -2.506749e-08, -1.539255e-08, -5.910174e-09, 
    5.910174e-09, 1.539255e-08, 2.506749e-08, 2.878978e-08, -7.008032e-09,
  7.008032e-09, -2.878978e-08, -2.506749e-08, -1.539255e-08, -5.910174e-09, 
    5.910174e-09, 1.539255e-08, 2.506749e-08, 2.878978e-08, -7.008032e-09,
  5.804671e-09, -2.381888e-08, -2.450905e-08, -1.50993e-08, -5.1423e-09, 
    5.1423e-09, 1.50993e-08, 2.450905e-08, 2.381888e-08, -5.804671e-09,
  0, -4.230289e-09, -1.879162e-08, -1.511646e-08, -4.975775e-09, 
    4.975775e-09, 1.511646e-08, 1.879162e-08, 4.230289e-09, 0,
  0, 2.319781e-09, -4.599584e-09, -4.862396e-09, -9.173195e-10, 9.173195e-10, 
    4.862396e-09, 4.599584e-09, -2.319781e-09, 0,
  0, 0, 0, 8.882792e-10, 2.049165e-10, -2.049165e-10, -8.882792e-10, 0, 0, 0,
  0, 0, 0, 4.980121e-05, 2.342554e-05, -2.342554e-05, -4.980121e-05, 0, 0, 0,
  0, -0.0001232052, 0.0005050731, -0.0001931989, -8.968446e-05, 8.968446e-05, 
    0.0001931989, -0.0005050731, 0.0001232052, 0,
  0, 0.0005791325, -0.002350952, -0.005442988, -0.001682935, 0.001682935, 
    0.005442988, 0.002350952, -0.0005791325, 0,
  0.0005110904, -0.0019067, -0.008924956, -0.004234629, -0.0008943132, 
    0.0008943132, 0.004234629, 0.008924956, 0.0019067, -0.0005110904,
  0.0009751136, -0.003646616, -0.009382538, -0.002442166, -0.0001501193, 
    0.0001501193, 0.002442166, 0.009382538, 0.003646616, -0.0009751136,
  0.0009751136, -0.003646616, -0.009382538, -0.002442166, -0.0001501193, 
    0.0001501193, 0.002442166, 0.009382538, 0.003646616, -0.0009751136,
  0.0005110904, -0.0019067, -0.008924956, -0.004234629, -0.0008943132, 
    0.0008943132, 0.004234629, 0.008924956, 0.0019067, -0.0005110904,
  0, 0.0005791325, -0.002350952, -0.005442988, -0.001682935, 0.001682935, 
    0.005442988, 0.002350952, -0.0005791325, 0,
  0, -0.0001232052, 0.0005050731, -0.0001931989, -8.968446e-05, 8.968446e-05, 
    0.0001931989, -0.0005050731, 0.0001232052, 0,
  0, 0, 0, 4.980121e-05, 2.342554e-05, -2.342554e-05, -4.980121e-05, 0, 0, 0,
  0, 0, 0, 4.618923e-05, 2.375904e-05, -2.375904e-05, -4.618923e-05, 0, 0, 0,
  0, -0.0001254825, 0.0005033801, -0.0001806051, -9.038047e-05, 9.038047e-05, 
    0.0001806051, -0.0005033801, 0.0001254825, 0,
  0, 0.0005774138, -0.002306366, -0.005381955, -0.001660131, 0.001660131, 
    0.005381955, 0.002306366, -0.0005774138, 0,
  0.0004972908, -0.001856323, -0.008823977, -0.004176188, -0.0008612028, 
    0.0008612028, 0.004176188, 0.008823977, 0.001856323, -0.0004972908,
  0.0009639504, -0.003599732, -0.009260577, -0.002364439, -0.0001416985, 
    0.0001416985, 0.002364439, 0.009260577, 0.003599732, -0.0009639504,
  0.0009639504, -0.003599732, -0.009260577, -0.002364439, -0.0001416985, 
    0.0001416985, 0.002364439, 0.009260577, 0.003599732, -0.0009639504,
  0.0004972908, -0.001856323, -0.008823977, -0.004176188, -0.0008612028, 
    0.0008612028, 0.004176188, 0.008823977, 0.001856323, -0.0004972908,
  0, 0.0005774138, -0.002306366, -0.005381955, -0.001660131, 0.001660131, 
    0.005381955, 0.002306366, -0.0005774138, 0,
  0, -0.0001254825, 0.0005033801, -0.0001806051, -9.038047e-05, 9.038047e-05, 
    0.0001806051, -0.0005033801, 0.0001254825, 0,
  0, 0, 0, 4.618923e-05, 2.375904e-05, -2.375904e-05, -4.618923e-05, 0, 0, 0,
  0, 0, 0, 4.035887e-05, 2.379059e-05, -2.379059e-05, -4.035887e-05, 0, 0, 0,
  0, -0.0001251925, 0.0004903096, -0.0001582718, -8.98889e-05, 8.98889e-05, 
    0.0001582718, -0.0004903096, 0.0001251925, 0,
  0, 0.0005597036, -0.002193888, -0.005192575, -0.001591897, 0.001591897, 
    0.005192575, 0.002193888, -0.0005597036, 0,
  0.0004646453, -0.001735174, -0.008513852, -0.0039785, -0.0007879224, 
    0.0007879224, 0.0039785, 0.008513852, 0.001735174, -0.0004646453,
  0.0009277874, -0.003462107, -0.008902945, -0.002171342, -0.0001243996, 
    0.0001243996, 0.002171342, 0.008902945, 0.003462107, -0.0009277874,
  0.0009277874, -0.003462107, -0.008902945, -0.002171342, -0.0001243996, 
    0.0001243996, 0.002171342, 0.008902945, 0.003462107, -0.0009277874,
  0.0004646453, -0.001735174, -0.008513852, -0.0039785, -0.0007879224, 
    0.0007879224, 0.0039785, 0.008513852, 0.001735174, -0.0004646453,
  0, 0.0005597036, -0.002193888, -0.005192575, -0.001591897, 0.001591897, 
    0.005192575, 0.002193888, -0.0005597036, 0,
  0, -0.0001251925, 0.0004903096, -0.0001582718, -8.98889e-05, 8.98889e-05, 
    0.0001582718, -0.0004903096, 0.0001251925, 0,
  0, 0, 0, 4.035887e-05, 2.379059e-05, -2.379059e-05, -4.035887e-05, 0, 0, 0,
  0, 0, 0, 3.402655e-05, 2.22479e-05, -2.22479e-05, -3.402655e-05, 0, 0, 0,
  0, -0.0001178382, 0.0004552921, -0.0001330857, -8.378804e-05, 8.378804e-05, 
    0.0001330857, -0.0004552921, 0.0001178382, 0,
  0, 0.0005156007, -0.001998015, -0.004806186, -0.001465671, 0.001465671, 
    0.004806186, 0.001998015, -0.0005156007, 0,
  0.0004163565, -0.001554788, -0.007881463, -0.003637122, -0.0006959632, 
    0.0006959632, 0.003637122, 0.007881463, 0.001554788, -0.0004163565,
  0.0008508377, -0.003174104, -0.008224366, -0.001920068, -0.0001036839, 
    0.0001036839, 0.001920068, 0.008224366, 0.003174104, -0.0008508377,
  0.0008508377, -0.003174104, -0.008224366, -0.001920068, -0.0001036839, 
    0.0001036839, 0.001920068, 0.008224366, 0.003174104, -0.0008508377,
  0.0004163565, -0.001554788, -0.007881463, -0.003637122, -0.0006959632, 
    0.0006959632, 0.003637122, 0.007881463, 0.001554788, -0.0004163565,
  0, 0.0005156007, -0.001998015, -0.004806186, -0.001465671, 0.001465671, 
    0.004806186, 0.001998015, -0.0005156007, 0,
  0, -0.0001178382, 0.0004552921, -0.0001330857, -8.378804e-05, 8.378804e-05, 
    0.0001330857, -0.0004552921, 0.0001178382, 0,
  0, 0, 0, 3.402655e-05, 2.22479e-05, -2.22479e-05, -3.402655e-05, 0, 0, 0,
  0, 0, 0, 2.754993e-05, 1.941581e-05, -1.941581e-05, -2.754993e-05, 0, 0, 0,
  0, -0.0001039136, 0.0003987052, -0.0001071937, -7.297657e-05, 7.297657e-05, 
    0.0001071937, -0.0003987052, 0.0001039136, 0,
  0, 0.000448019, -0.001725244, -0.004214888, -0.001280167, 0.001280167, 
    0.004214888, 0.001725244, -0.000448019, 0,
  0.000355047, -0.001325687, -0.006912369, -0.003158372, -0.000590838, 
    0.000590838, 0.003158372, 0.006912369, 0.001325687, -0.000355047,
  0.0007369739, -0.002749153, -0.007209442, -0.001628536, -8.356683e-05, 
    8.356683e-05, 0.001628536, 0.007209442, 0.002749153, -0.0007369739,
  0.0007369739, -0.002749153, -0.007209442, -0.001628536, -8.356683e-05, 
    8.356683e-05, 0.001628536, 0.007209442, 0.002749153, -0.0007369739,
  0.000355047, -0.001325687, -0.006912369, -0.003158372, -0.000590838, 
    0.000590838, 0.003158372, 0.006912369, 0.001325687, -0.000355047,
  0, 0.000448019, -0.001725244, -0.004214888, -0.001280167, 0.001280167, 
    0.004214888, 0.001725244, -0.000448019, 0,
  0, -0.0001039136, 0.0003987052, -0.0001071937, -7.297657e-05, 7.297657e-05, 
    0.0001071937, -0.0003987052, 0.0001039136, 0,
  0, 0, 0, 2.754993e-05, 1.941581e-05, -1.941581e-05, -2.754993e-05, 0, 0, 0,
  0, 0, 0, 2.118585e-05, 1.583643e-05, -1.583643e-05, -2.118585e-05, 0, 0, 0,
  0, -8.559917e-05, 0.000327143, -8.191521e-05, -5.942961e-05, 5.942961e-05, 
    8.191521e-05, -0.000327143, 8.559917e-05, 0,
  0, 0.0003653085, -0.001401504, -0.00347171, -0.001050762, 0.001050762, 
    0.00347171, 0.001401504, -0.0003653085, 0,
  0.0002855763, -0.001066172, -0.005693769, -0.002579907, -0.0004757417, 
    0.0004757417, 0.002579907, 0.005693769, 0.001066172, -0.0002855763,
  0.0005992496, -0.002235452, -0.005938564, -0.001308785, -6.508073e-05, 
    6.508073e-05, 0.001308785, 0.005938564, 0.002235452, -0.0005992496,
  0.0005992496, -0.002235452, -0.005938564, -0.001308785, -6.508073e-05, 
    6.508073e-05, 0.001308785, 0.005938564, 0.002235452, -0.0005992496,
  0.0002855763, -0.001066172, -0.005693769, -0.002579907, -0.0004757417, 
    0.0004757417, 0.002579907, 0.005693769, 0.001066172, -0.0002855763,
  0, 0.0003653085, -0.001401504, -0.00347171, -0.001050762, 0.001050762, 
    0.00347171, 0.001401504, -0.0003653085, 0,
  0, -8.559917e-05, 0.000327143, -8.191521e-05, -5.942961e-05, 5.942961e-05, 
    8.191521e-05, -0.000327143, 8.559917e-05, 0,
  0, 0, 0, 2.118585e-05, 1.583643e-05, -1.583643e-05, -2.118585e-05, 0, 0, 0,
  0, 0, 0, 1.51612e-05, 1.189718e-05, -1.189718e-05, -1.51612e-05, 0, 0, 0,
  0, -6.485327e-05, 0.0002472673, -5.821702e-05, -4.458491e-05, 4.458491e-05, 
    5.821702e-05, -0.0002472673, 6.485327e-05, 0,
  0, 0.0002748477, -0.00105202, -0.0026385, -0.000795964, 0.000795964, 
    0.0026385, 0.00105202, -0.0002748477, 0,
  0.00021265, -0.0007938269, -0.004327347, -0.001945966, -0.0003554224, 
    0.0003554224, 0.001945966, 0.004327347, 0.0007938269, -0.00021265,
  0.000449594, -0.001677288, -0.004513612, -0.0009755426, -4.778522e-05, 
    4.778522e-05, 0.0009755426, 0.004513612, 0.001677288, -0.000449594,
  0.000449594, -0.001677288, -0.004513612, -0.0009755426, -4.778522e-05, 
    4.778522e-05, 0.0009755426, 0.004513612, 0.001677288, -0.000449594,
  0.00021265, -0.0007938269, -0.004327347, -0.001945966, -0.0003554224, 
    0.0003554224, 0.001945966, 0.004327347, 0.0007938269, -0.00021265,
  0, 0.0002748477, -0.00105202, -0.0026385, -0.000795964, 0.000795964, 
    0.0026385, 0.00105202, -0.0002748477, 0,
  0, -6.485327e-05, 0.0002472673, -5.821702e-05, -4.458491e-05, 4.458491e-05, 
    5.821702e-05, -0.0002472673, 6.485327e-05, 0,
  0, 0, 0, 1.51612e-05, 1.189718e-05, -1.189718e-05, -1.51612e-05, 0, 0, 0,
  0, 0, 0, 9.574579e-06, 7.856769e-06, -7.856769e-06, -9.574579e-06, 0, 0, 0,
  0, -4.311253e-05, 0.0001641228, -3.649069e-05, -2.940429e-05, 2.940429e-05, 
    3.649069e-05, -0.0001641228, 4.311253e-05, 0,
  0, 0.0001818528, -0.0006950366, -0.001764653, -0.0005308443, 0.0005308443, 
    0.001764653, 0.0006950366, -0.0001818528, 0,
  0.0001395506, -0.000520897, -0.002894199, -0.001292788, -0.0002344245, 
    0.0002344245, 0.001292788, 0.002894199, 0.000520897, -0.0001395506,
  0.0002966736, -0.001106895, -0.003019516, -0.0006419583, -3.13057e-05, 
    3.13057e-05, 0.0006419583, 0.003019516, 0.001106895, -0.0002966736,
  0.0002966736, -0.001106895, -0.003019516, -0.0006419583, -3.13057e-05, 
    3.13057e-05, 0.0006419583, 0.003019516, 0.001106895, -0.0002966736,
  0.0001395506, -0.000520897, -0.002894199, -0.001292788, -0.0002344245, 
    0.0002344245, 0.001292788, 0.002894199, 0.000520897, -0.0001395506,
  0, 0.0001818528, -0.0006950366, -0.001764653, -0.0005308443, 0.0005308443, 
    0.001764653, 0.0006950366, -0.0001818528, 0,
  0, -4.311253e-05, 0.0001641228, -3.649069e-05, -2.940429e-05, 2.940429e-05, 
    3.649069e-05, -0.0001641228, 4.311253e-05, 0,
  0, 0, 0, 9.574579e-06, 7.856769e-06, -7.856769e-06, -9.574579e-06, 0, 0, 0,
  0, 0, 0, 4.472497e-06, 3.866233e-06, -3.866233e-06, -4.472497e-06, 0, 0, 0,
  0, -2.130998e-05, 8.10249e-05, -1.689914e-05, -1.444882e-05, 1.444882e-05, 
    1.689914e-05, -8.10249e-05, 2.130998e-05, 0,
  0, 8.958419e-05, -0.0003420194, -0.0008810312, -0.0002647389, 0.0002647389, 
    0.0008810312, 0.0003420194, -8.958419e-05, 0,
  6.823079e-05, -0.0002546627, -0.001444988, -0.0006430848, -0.0001158388, 
    0.0001158388, 0.0006430848, 0.001444988, 0.0002546627, -6.823079e-05,
  0.0001458607, -0.0005442753, -0.001509905, -0.000316673, -1.546205e-05, 
    1.546205e-05, 0.000316673, 0.001509905, 0.0005442753, -0.0001458607,
  0.0001458607, -0.0005442753, -0.001509905, -0.000316673, -1.546205e-05, 
    1.546205e-05, 0.000316673, 0.001509905, 0.0005442753, -0.0001458607,
  6.823079e-05, -0.0002546627, -0.001444988, -0.0006430848, -0.0001158388, 
    0.0001158388, 0.0006430848, 0.001444988, 0.0002546627, -6.823079e-05,
  0, 8.958419e-05, -0.0003420194, -0.0008810312, -0.0002647389, 0.0002647389, 
    0.0008810312, 0.0003420194, -8.958419e-05, 0,
  0, -2.130998e-05, 8.10249e-05, -1.689914e-05, -1.444882e-05, 1.444882e-05, 
    1.689914e-05, -8.10249e-05, 2.130998e-05, 0,
  0, 0, 0, 4.472497e-06, 3.866233e-06, -3.866233e-06, -4.472497e-06, 0, 0, 0,
  0, 0, 0, 8.882624e-10, 2.051505e-10, -2.051505e-10, -8.882624e-10, 0, 0, 0,
  0, 2.323635e-09, -4.609836e-09, -4.868089e-09, -9.183869e-10, 9.183869e-10, 
    4.868089e-09, 4.609836e-09, -2.323635e-09, 0,
  0, -4.243433e-09, -1.879897e-08, -1.509725e-08, -4.972821e-09, 
    4.972821e-09, 1.509725e-08, 1.879897e-08, 4.243433e-09, 0,
  5.808406e-09, -2.384734e-08, -2.446902e-08, -1.507616e-08, -5.141223e-09, 
    5.141223e-09, 1.507616e-08, 2.446902e-08, 2.384734e-08, -5.808406e-09,
  7.008185e-09, -2.881204e-08, -2.500002e-08, -1.539884e-08, -5.929314e-09, 
    5.929314e-09, 1.539884e-08, 2.500002e-08, 2.881204e-08, -7.008185e-09,
  7.008185e-09, -2.881204e-08, -2.500002e-08, -1.539884e-08, -5.929314e-09, 
    5.929314e-09, 1.539884e-08, 2.500002e-08, 2.881204e-08, -7.008185e-09,
  5.808406e-09, -2.384734e-08, -2.446902e-08, -1.507616e-08, -5.141223e-09, 
    5.141223e-09, 1.507616e-08, 2.446902e-08, 2.384734e-08, -5.808406e-09,
  0, -4.243433e-09, -1.879897e-08, -1.509725e-08, -4.972821e-09, 
    4.972821e-09, 1.509725e-08, 1.879897e-08, 4.243433e-09, 0,
  0, 2.323635e-09, -4.609836e-09, -4.868089e-09, -9.183869e-10, 9.183869e-10, 
    4.868089e-09, 4.609836e-09, -2.323635e-09, 0,
  0, 0, 0, 8.882624e-10, 2.051505e-10, -2.051505e-10, -8.882624e-10, 0, 0, 0 ;

 velnorm =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0008830973, 0.01197786, 0.05273421, 0.05273421, 0.01197786, 
    0.0008830973, 0, 0,
  0, 0.0008830973, 0.01182386, 0.01156157, 0.01126752, 0.01126752, 
    0.01156157, 0.01182386, 0.0008830973, 0,
  0, 0.01197786, 0.01156157, 0.006455652, 0.002303052, 0.002303052, 
    0.006455652, 0.01156157, 0.01197786, 0,
  0, 0.05273421, 0.01126752, 0.002303052, 0.0002353543, 0.0002353543, 
    0.002303052, 0.01126752, 0.05273421, 0,
  0, 0.05273421, 0.01126752, 0.002303052, 0.0002353543, 0.0002353543, 
    0.002303052, 0.01126752, 0.05273421, 0,
  0, 0.01197786, 0.01156157, 0.006455652, 0.002303052, 0.002303052, 
    0.006455652, 0.01156157, 0.01197786, 0,
  0, 0.0008830973, 0.01182386, 0.01156157, 0.01126752, 0.01126752, 
    0.01156157, 0.01182386, 0.0008830973, 0,
  0, 0, 0.0008830973, 0.01197786, 0.05273421, 0.05273421, 0.01197786, 
    0.0008830973, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0009323089, 0.01184183, 0.05202222, 0.05202222, 0.01184183, 
    0.0009323089, 0, 0,
  0, 0.0009323089, 0.01171938, 0.01147223, 0.01100237, 0.01100237, 
    0.01147223, 0.01171938, 0.0009323089, 0,
  0, 0.01184183, 0.01147223, 0.006322624, 0.002244861, 0.002244861, 
    0.006322624, 0.01147223, 0.01184183, 0,
  0, 0.05202222, 0.01100237, 0.002244861, 0.0002181856, 0.0002181856, 
    0.002244861, 0.01100237, 0.05202222, 0,
  0, 0.05202222, 0.01100237, 0.002244861, 0.0002181856, 0.0002181856, 
    0.002244861, 0.01100237, 0.05202222, 0,
  0, 0.01184183, 0.01147223, 0.006322624, 0.002244861, 0.002244861, 
    0.006322624, 0.01147223, 0.01184183, 0,
  0, 0.0009323089, 0.01171938, 0.01147223, 0.01100237, 0.01100237, 
    0.01147223, 0.01171938, 0.0009323089, 0,
  0, 0, 0.0009323089, 0.01184183, 0.05202222, 0.05202222, 0.01184183, 
    0.0009323089, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.001014795, 0.01139397, 0.04994358, 0.04994358, 0.01139397, 
    0.001014795, 0, 0,
  0, 0.001014795, 0.01133603, 0.01110497, 0.0102722, 0.0102722, 0.01110497, 
    0.01133603, 0.001014795, 0,
  0, 0.01139397, 0.01110497, 0.005966518, 0.002096084, 0.002096084, 
    0.005966518, 0.01110497, 0.01139397, 0,
  0, 0.04994358, 0.0102722, 0.002096084, 0.0001827411, 0.0001827411, 
    0.002096084, 0.0102722, 0.04994358, 0,
  0, 0.04994358, 0.0102722, 0.002096084, 0.0001827411, 0.0001827411, 
    0.002096084, 0.0102722, 0.04994358, 0,
  0, 0.01139397, 0.01110497, 0.005966518, 0.002096084, 0.002096084, 
    0.005966518, 0.01110497, 0.01139397, 0,
  0, 0.001014795, 0.01133603, 0.01110497, 0.0102722, 0.0102722, 0.01110497, 
    0.01133603, 0.001014795, 0,
  0, 0, 0.001014795, 0.01139397, 0.04994358, 0.04994358, 0.01139397, 
    0.001014795, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.001033265, 0.01046101, 0.04609964, 0.04609964, 0.01046101, 
    0.001033265, 0, 0,
  0, 0.001033265, 0.01047179, 0.01027817, 0.009208306, 0.009208306, 
    0.01027817, 0.01047179, 0.001033265, 0,
  0, 0.01046101, 0.01027817, 0.005417457, 0.001884199, 0.001884199, 
    0.005417457, 0.01027817, 0.01046101, 0,
  0, 0.04609964, 0.009208306, 0.001884199, 0.0001447224, 0.0001447224, 
    0.001884199, 0.009208306, 0.04609964, 0,
  0, 0.04609964, 0.009208306, 0.001884199, 0.0001447224, 0.0001447224, 
    0.001884199, 0.009208306, 0.04609964, 0,
  0, 0.01046101, 0.01027817, 0.005417457, 0.001884199, 0.001884199, 
    0.005417457, 0.01027817, 0.01046101, 0,
  0, 0.001033265, 0.01047179, 0.01027817, 0.009208306, 0.009208306, 
    0.01027817, 0.01047179, 0.001033265, 0,
  0, 0, 0.001033265, 0.01046101, 0.04609964, 0.04609964, 0.01046101, 
    0.001033265, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0009653685, 0.009075353, 0.04037431, 0.04037431, 0.009075353, 
    0.0009653685, 0, 0,
  0, 0.0009653685, 0.009144534, 0.008990949, 0.007871899, 0.007871899, 
    0.008990949, 0.009144534, 0.0009653685, 0,
  0, 0.009075353, 0.008990949, 0.004682323, 0.001620586, 0.001620586, 
    0.004682323, 0.008990949, 0.009075353, 0,
  0, 0.04037431, 0.007871899, 0.001620586, 0.0001110042, 0.0001110042, 
    0.001620586, 0.007871899, 0.04037431, 0,
  0, 0.04037431, 0.007871899, 0.001620586, 0.0001110042, 0.0001110042, 
    0.001620586, 0.007871899, 0.04037431, 0,
  0, 0.009075353, 0.008990949, 0.004682323, 0.001620586, 0.001620586, 
    0.004682323, 0.008990949, 0.009075353, 0,
  0, 0.0009653685, 0.009144534, 0.008990949, 0.007871899, 0.007871899, 
    0.008990949, 0.009144534, 0.0009653685, 0,
  0, 0, 0.0009653685, 0.009075353, 0.04037431, 0.04037431, 0.009075353, 
    0.0009653685, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0008303312, 0.007388042, 0.03320354, 0.03320354, 0.007388042, 
    0.0008303312, 0, 0,
  0, 0.0008303312, 0.007490865, 0.007374792, 0.006346367, 0.006346367, 
    0.007374792, 0.007490865, 0.0008303312, 0,
  0, 0.007388042, 0.007374792, 0.003809904, 0.001317447, 0.001317447, 
    0.003809904, 0.007374792, 0.007388042, 0,
  0, 0.03320354, 0.006346367, 0.001317447, 8.250551e-05, 8.250551e-05, 
    0.001317447, 0.006346367, 0.03320354, 0,
  0, 0.03320354, 0.006346367, 0.001317447, 8.250551e-05, 8.250551e-05, 
    0.001317447, 0.006346367, 0.03320354, 0,
  0, 0.007388042, 0.007374792, 0.003809904, 0.001317447, 0.001317447, 
    0.003809904, 0.007374792, 0.007388042, 0,
  0, 0.0008303312, 0.007490865, 0.007374792, 0.006346367, 0.006346367, 
    0.007374792, 0.007490865, 0.0008303312, 0,
  0, 0, 0.0008303312, 0.007388042, 0.03320354, 0.03320354, 0.007388042, 
    0.0008303312, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0006501422, 0.005544633, 0.02515636, 0.02515636, 0.005544633, 
    0.0006501422, 0, 0,
  0, 0.0006501422, 0.005653069, 0.005571141, 0.004729439, 0.004729439, 
    0.005571141, 0.005653069, 0.0006501422, 0,
  0, 0.005544633, 0.005571141, 0.002861537, 0.000990534, 0.000990534, 
    0.002861537, 0.005571141, 0.005544633, 0,
  0, 0.02515636, 0.004729439, 0.000990534, 5.801751e-05, 5.801751e-05, 
    0.000990534, 0.004729439, 0.02515636, 0,
  0, 0.02515636, 0.004729439, 0.000990534, 5.801751e-05, 5.801751e-05, 
    0.000990534, 0.004729439, 0.02515636, 0,
  0, 0.005544633, 0.005571141, 0.002861537, 0.000990534, 0.000990534, 
    0.002861537, 0.005571141, 0.005544633, 0,
  0, 0.0006501422, 0.005653069, 0.005571141, 0.004729439, 0.004729439, 
    0.005571141, 0.005653069, 0.0006501422, 0,
  0, 0, 0.0006501422, 0.005544633, 0.02515636, 0.02515636, 0.005544633, 
    0.0006501422, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0004431279, 0.003654536, 0.01672114, 0.01672114, 0.003654536, 
    0.0004431279, 0, 0,
  0, 0.0004431279, 0.003743982, 0.003692668, 0.003100349, 0.003100349, 
    0.003692668, 0.003743982, 0.0004431279, 0,
  0, 0.003654536, 0.003692668, 0.001888427, 0.0006548685, 0.0006548685, 
    0.001888427, 0.003692668, 0.003654536, 0,
  0, 0.01672114, 0.003100349, 0.0006548685, 3.647256e-05, 3.647256e-05, 
    0.0006548685, 0.003100349, 0.01672114, 0,
  0, 0.01672114, 0.003100349, 0.0006548685, 3.647256e-05, 3.647256e-05, 
    0.0006548685, 0.003100349, 0.01672114, 0,
  0, 0.003654536, 0.003692668, 0.001888427, 0.0006548685, 0.0006548685, 
    0.001888427, 0.003692668, 0.003654536, 0,
  0, 0.0004431279, 0.003743982, 0.003692668, 0.003100349, 0.003100349, 
    0.003692668, 0.003743982, 0.0004431279, 0,
  0, 0, 0.0004431279, 0.003654536, 0.01672114, 0.01672114, 0.003654536, 
    0.0004431279, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0002231378, 0.001791215, 0.008255952, 0.008255952, 0.001791215, 
    0.0002231378, 0, 0,
  0, 0.0002231378, 0.001842662, 0.001818561, 0.00151299, 0.00151299, 
    0.001818561, 0.001842662, 0.0002231378, 0,
  0, 0.001791215, 0.001818561, 0.0009268459, 0.0003220633, 0.0003220633, 
    0.0009268459, 0.001818561, 0.001791215, 0,
  0, 0.008255952, 0.00151299, 0.0003220633, 1.725464e-05, 1.725464e-05, 
    0.0003220633, 0.00151299, 0.008255952, 0,
  0, 0.008255952, 0.00151299, 0.0003220633, 1.725464e-05, 1.725464e-05, 
    0.0003220633, 0.00151299, 0.008255952, 0,
  0, 0.001791215, 0.001818561, 0.0009268459, 0.0003220633, 0.0003220633, 
    0.0009268459, 0.001818561, 0.001791215, 0,
  0, 0.0002231378, 0.001842662, 0.001818561, 0.00151299, 0.00151299, 
    0.001818561, 0.001842662, 0.0002231378, 0,
  0, 0, 0.0002231378, 0.001791215, 0.008255952, 0.008255952, 0.001791215, 
    0.0002231378, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.71268e-08, 3.457684e-08, 5.11253e-08, 5.11253e-08, 3.457684e-08, 
    1.71268e-08, 0, 0,
  0, 1.71268e-08, 3.330913e-08, 2.944244e-08, 2.770732e-08, 2.770732e-08, 
    2.944244e-08, 3.330913e-08, 1.71268e-08, 0,
  0, 3.457684e-08, 2.944244e-08, 2.202386e-08, 1.566339e-08, 1.566339e-08, 
    2.202386e-08, 2.944244e-08, 3.457684e-08, 0,
  0, 5.11253e-08, 2.770732e-08, 1.566339e-08, 8.286722e-09, 8.286722e-09, 
    1.566339e-08, 2.770732e-08, 5.11253e-08, 0,
  0, 5.11253e-08, 2.770732e-08, 1.566339e-08, 8.286722e-09, 8.286722e-09, 
    1.566339e-08, 2.770732e-08, 5.11253e-08, 0,
  0, 3.457684e-08, 2.944244e-08, 2.202386e-08, 1.566339e-08, 1.566339e-08, 
    2.202386e-08, 2.944244e-08, 3.457684e-08, 0,
  0, 1.71268e-08, 3.330913e-08, 2.944244e-08, 2.770732e-08, 2.770732e-08, 
    2.944244e-08, 3.330913e-08, 1.71268e-08, 0,
  0, 0, 1.71268e-08, 3.457684e-08, 5.11253e-08, 5.11253e-08, 3.457684e-08, 
    1.71268e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002908382, 0.002908382, 0, 0, 0, 0,
  0, 0, 0.001654083, 0.01411019, 0.01095244, 0.01095244, 0.01411019, 
    0.001654083, 0, 0,
  0, 0.001654083, 0.01179826, 0.01155781, 0.01098661, 0.01098661, 0.01155781, 
    0.01179826, 0.001654083, 0,
  0, 0.01411019, 0.01155781, 0.006386738, 0.00244144, 0.00244144, 
    0.006386738, 0.01155781, 0.01411019, 0,
  0.002908382, 0.01095244, 0.01098661, 0.00244144, 0.0001921582, 
    0.0001921582, 0.00244144, 0.01098661, 0.01095244, 0.002908382,
  0.002908382, 0.01095244, 0.01098661, 0.00244144, 0.0001921582, 
    0.0001921582, 0.00244144, 0.01098661, 0.01095244, 0.002908382,
  0, 0.01411019, 0.01155781, 0.006386738, 0.00244144, 0.00244144, 
    0.006386738, 0.01155781, 0.01411019, 0,
  0, 0.001654083, 0.01179826, 0.01155781, 0.01098661, 0.01098661, 0.01155781, 
    0.01179826, 0.001654083, 0,
  0, 0, 0.001654083, 0.01411019, 0.01095244, 0.01095244, 0.01411019, 
    0.001654083, 0, 0,
  0, 0, 0, 0, 0.002908382, 0.002908382, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002903924, 0.002903924, 0, 0, 0, 0,
  0, 0, 0.001731203, 0.01401759, 0.01088206, 0.01088206, 0.01401759, 
    0.001731203, 0, 0,
  0, 0.001731203, 0.01170186, 0.01145189, 0.01087959, 0.01087959, 0.01145189, 
    0.01170186, 0.001731203, 0,
  0, 0.01401759, 0.01145189, 0.006260482, 0.002352321, 0.002352321, 
    0.006260482, 0.01145189, 0.01401759, 0,
  0.002903924, 0.01088206, 0.01087959, 0.002352321, 0.0001844815, 
    0.0001844815, 0.002352321, 0.01087959, 0.01088206, 0.002903924,
  0.002903924, 0.01088206, 0.01087959, 0.002352321, 0.0001844815, 
    0.0001844815, 0.002352321, 0.01087959, 0.01088206, 0.002903924,
  0, 0.01401759, 0.01145189, 0.006260482, 0.002352321, 0.002352321, 
    0.006260482, 0.01145189, 0.01401759, 0,
  0, 0.001731203, 0.01170186, 0.01145189, 0.01087959, 0.01087959, 0.01145189, 
    0.01170186, 0.001731203, 0,
  0, 0, 0.001731203, 0.01401759, 0.01088206, 0.01088206, 0.01401759, 
    0.001731203, 0, 0,
  0, 0, 0, 0, 0.002903924, 0.002903924, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002813153, 0.002813153, 0, 0, 0, 0,
  0, 0, 0.001828402, 0.01359599, 0.01051697, 0.01051697, 0.01359599, 
    0.001828402, 0, 0,
  0, 0.001828402, 0.01133093, 0.01105687, 0.01044887, 0.01044887, 0.01105687, 
    0.01133093, 0.001828402, 0,
  0, 0.01359599, 0.01105687, 0.00591659, 0.002146706, 0.002146706, 
    0.00591659, 0.01105687, 0.01359599, 0,
  0.002813153, 0.01051697, 0.01044887, 0.002146706, 0.0001649879, 
    0.0001649879, 0.002146706, 0.01044887, 0.01051697, 0.002813153,
  0.002813153, 0.01051697, 0.01044887, 0.002146706, 0.0001649879, 
    0.0001649879, 0.002146706, 0.01044887, 0.01051697, 0.002813153,
  0, 0.01359599, 0.01105687, 0.00591659, 0.002146706, 0.002146706, 
    0.00591659, 0.01105687, 0.01359599, 0,
  0, 0.001828402, 0.01133093, 0.01105687, 0.01044887, 0.01044887, 0.01105687, 
    0.01133093, 0.001828402, 0,
  0, 0, 0.001828402, 0.01359599, 0.01051697, 0.01051697, 0.01359599, 
    0.001828402, 0, 0,
  0, 0, 0, 0, 0.002813153, 0.002813153, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002594745, 0.002594745, 0, 0, 0, 0,
  0, 0, 0.001811954, 0.01257066, 0.009690557, 0.009690557, 0.01257066, 
    0.001811954, 0, 0,
  0, 0.001811954, 0.01048287, 0.01020302, 0.009611952, 0.009611952, 
    0.01020302, 0.01048287, 0.001811954, 0,
  0, 0.01257066, 0.01020302, 0.005382852, 0.001889069, 0.001889069, 
    0.005382852, 0.01020302, 0.01257066, 0,
  0.002594745, 0.009690557, 0.009611952, 0.001889069, 0.0001393725, 
    0.0001393725, 0.001889069, 0.009611952, 0.009690557, 0.002594745,
  0.002594745, 0.009690557, 0.009611952, 0.001889069, 0.0001393725, 
    0.0001393725, 0.001889069, 0.009611952, 0.009690557, 0.002594745,
  0, 0.01257066, 0.01020302, 0.005382852, 0.001889069, 0.001889069, 
    0.005382852, 0.01020302, 0.01257066, 0,
  0, 0.001811954, 0.01048287, 0.01020302, 0.009611952, 0.009611952, 
    0.01020302, 0.01048287, 0.001811954, 0,
  0, 0, 0.001811954, 0.01257066, 0.009690557, 0.009690557, 0.01257066, 
    0.001811954, 0, 0,
  0, 0, 0, 0, 0.002594745, 0.002594745, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002259675, 0.002259675, 0, 0, 0, 0,
  0, 0, 0.001664985, 0.01097924, 0.008435003, 0.008435003, 0.01097924, 
    0.001664985, 0, 0,
  0, 0.001664985, 0.009167681, 0.008902882, 0.008383372, 0.008383372, 
    0.008902882, 0.009167681, 0.001664985, 0,
  0, 0.01097924, 0.008902882, 0.004660707, 0.001597729, 0.001597729, 
    0.004660707, 0.008902882, 0.01097924, 0,
  0.002259675, 0.008435003, 0.008383372, 0.001597729, 0.0001130466, 
    0.0001130466, 0.001597729, 0.008383372, 0.008435003, 0.002259675,
  0.002259675, 0.008435003, 0.008383372, 0.001597729, 0.0001130466, 
    0.0001130466, 0.001597729, 0.008383372, 0.008435003, 0.002259675,
  0, 0.01097924, 0.008902882, 0.004660707, 0.001597729, 0.001597729, 
    0.004660707, 0.008902882, 0.01097924, 0,
  0, 0.001664985, 0.009167681, 0.008902882, 0.008383372, 0.008383372, 
    0.008902882, 0.009167681, 0.001664985, 0,
  0, 0, 0.001664985, 0.01097924, 0.008435003, 0.008435003, 0.01097924, 
    0.001664985, 0, 0,
  0, 0, 0, 0, 0.002259675, 0.002259675, 0, 0, 0, 0,
  0, 0, 0, 0, 0.001845607, 0.001845607, 0, 0, 0, 0,
  0, 0, 0.001416923, 0.00899412, 0.006887729, 0.006887729, 0.00899412, 
    0.001416923, 0, 0,
  0, 0.001416923, 0.007520497, 0.007288414, 0.006868142, 0.006868142, 
    0.007288414, 0.007520497, 0.001416923, 0,
  0, 0.00899412, 0.007288414, 0.003798154, 0.00128172, 0.00128172, 
    0.003798154, 0.007288414, 0.00899412, 0,
  0.001845607, 0.006887729, 0.006868142, 0.00128172, 8.812103e-05, 
    8.812103e-05, 0.00128172, 0.006868142, 0.006887729, 0.001845607,
  0.001845607, 0.006887729, 0.006868142, 0.00128172, 8.812103e-05, 
    8.812103e-05, 0.00128172, 0.006868142, 0.006887729, 0.001845607,
  0, 0.00899412, 0.007288414, 0.003798154, 0.00128172, 0.00128172, 
    0.003798154, 0.007288414, 0.00899412, 0,
  0, 0.001416923, 0.007520497, 0.007288414, 0.006868142, 0.006868142, 
    0.007288414, 0.007520497, 0.001416923, 0,
  0, 0, 0.001416923, 0.00899412, 0.006887729, 0.006887729, 0.00899412, 
    0.001416923, 0, 0,
  0, 0, 0, 0, 0.001845607, 0.001845607, 0, 0, 0, 0,
  0, 0, 0, 0, 0.00138911, 0.00138911, 0, 0, 0, 0,
  0, 0, 0.001101479, 0.00678921, 0.005183605, 0.005183605, 0.00678921, 
    0.001101479, 0, 0,
  0, 0.001101479, 0.005684117, 0.005498307, 0.005187146, 0.005187146, 
    0.005498307, 0.005684117, 0.001101479, 0,
  0, 0.00678921, 0.005498307, 0.002856744, 0.000953436, 0.000953436, 
    0.002856744, 0.005498307, 0.00678921, 0,
  0.00138911, 0.005183605, 0.005187146, 0.000953436, 6.451798e-05, 
    6.451798e-05, 0.000953436, 0.005187146, 0.005183605, 0.00138911,
  0.00138911, 0.005183605, 0.005187146, 0.000953436, 6.451798e-05, 
    6.451798e-05, 0.000953436, 0.005187146, 0.005183605, 0.00138911,
  0, 0.00678921, 0.005498307, 0.002856744, 0.000953436, 0.000953436, 
    0.002856744, 0.005498307, 0.00678921, 0,
  0, 0.001101479, 0.005684117, 0.005498307, 0.005187146, 0.005187146, 
    0.005498307, 0.005684117, 0.001101479, 0,
  0, 0, 0.001101479, 0.00678921, 0.005183605, 0.005183605, 0.00678921, 
    0.001101479, 0, 0,
  0, 0, 0, 0, 0.00138911, 0.00138911, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0009180843, 0.0009180843, 0, 0, 0, 0,
  0, 0, 0.0007471829, 0.004500463, 0.003425877, 0.003425877, 0.004500463, 
    0.0007471829, 0, 0,
  0, 0.0007471829, 0.003772113, 0.003642041, 0.003440066, 0.003440066, 
    0.003642041, 0.003772113, 0.0007471829, 0,
  0, 0.004500463, 0.003642041, 0.001888091, 0.0006249872, 0.0006249872, 
    0.001888091, 0.003642041, 0.004500463, 0,
  0.0009180843, 0.003425877, 0.003440066, 0.0006249872, 4.197975e-05, 
    4.197975e-05, 0.0006249872, 0.003440066, 0.003425877, 0.0009180843,
  0.0009180843, 0.003425877, 0.003440066, 0.0006249872, 4.197975e-05, 
    4.197975e-05, 0.0006249872, 0.003440066, 0.003425877, 0.0009180843,
  0, 0.004500463, 0.003642041, 0.001888091, 0.0006249872, 0.0006249872, 
    0.001888091, 0.003642041, 0.004500463, 0,
  0, 0.0007471829, 0.003772113, 0.003642041, 0.003440066, 0.003440066, 
    0.003642041, 0.003772113, 0.0007471829, 0,
  0, 0, 0.0007471829, 0.004500463, 0.003425877, 0.003425877, 0.004500463, 
    0.0007471829, 0, 0,
  0, 0, 0, 0, 0.0009180843, 0.0009180843, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0004514559, 0.0004514559, 0, 0, 0, 0,
  0, 0, 0.0003755426, 0.002220839, 0.001684703, 0.001684703, 0.002220839, 
    0.0003755426, 0, 0,
  0, 0.0003755426, 0.00186301, 0.001795301, 0.00169777, 0.00169777, 
    0.001795301, 0.00186301, 0.0003755426, 0,
  0, 0.002220839, 0.001795301, 0.0009289205, 0.00030548, 0.00030548, 
    0.0009289205, 0.001795301, 0.002220839, 0,
  0.0004514559, 0.001684703, 0.00169777, 0.00030548, 2.047736e-05, 
    2.047736e-05, 0.00030548, 0.00169777, 0.001684703, 0.0004514559,
  0.0004514559, 0.001684703, 0.00169777, 0.00030548, 2.047736e-05, 
    2.047736e-05, 0.00030548, 0.00169777, 0.001684703, 0.0004514559,
  0, 0.002220839, 0.001795301, 0.0009289205, 0.00030548, 0.00030548, 
    0.0009289205, 0.001795301, 0.002220839, 0,
  0, 0.0003755426, 0.00186301, 0.001795301, 0.00169777, 0.00169777, 
    0.001795301, 0.00186301, 0.0003755426, 0,
  0, 0, 0.0003755426, 0.002220839, 0.001684703, 0.001684703, 0.002220839, 
    0.0003755426, 0, 0,
  0, 0, 0, 0, 0.0004514559, 0.0004514559, 0, 0, 0, 0,
  0, 0, 0, 0, 8.245442e-09, 8.245442e-09, 0, 0, 0, 0,
  0, 0, 1.727301e-08, 3.455769e-08, 3.656173e-08, 3.656173e-08, 3.455769e-08, 
    1.727301e-08, 0, 0,
  0, 1.727301e-08, 3.314176e-08, 2.963724e-08, 2.649972e-08, 2.649972e-08, 
    2.963724e-08, 3.314176e-08, 1.727301e-08, 0,
  0, 3.455769e-08, 2.963724e-08, 2.184066e-08, 1.610376e-08, 1.610376e-08, 
    2.184066e-08, 2.963724e-08, 3.455769e-08, 0,
  8.245442e-09, 3.656173e-08, 2.649972e-08, 1.610376e-08, 8.079599e-09, 
    8.079599e-09, 1.610376e-08, 2.649972e-08, 3.656173e-08, 8.245442e-09,
  8.245442e-09, 3.656173e-08, 2.649972e-08, 1.610376e-08, 8.079599e-09, 
    8.079599e-09, 1.610376e-08, 2.649972e-08, 3.656173e-08, 8.245442e-09,
  0, 3.455769e-08, 2.963724e-08, 2.184066e-08, 1.610376e-08, 1.610376e-08, 
    2.184066e-08, 2.963724e-08, 3.455769e-08, 0,
  0, 1.727301e-08, 3.314176e-08, 2.963724e-08, 2.649972e-08, 2.649972e-08, 
    2.963724e-08, 3.314176e-08, 1.727301e-08, 0,
  0, 0, 1.727301e-08, 3.455769e-08, 3.656173e-08, 3.656173e-08, 3.455769e-08, 
    1.727301e-08, 0, 0,
  0, 0, 0, 0, 8.245442e-09, 8.245442e-09, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002910513, 0.002910513, 0, 0, 0, 0,
  0, 0, 0.001642336, 0.01412936, 0.01096149, 0.01096149, 0.01412936, 
    0.001642336, 0, 0,
  0, 0.001642336, 0.01180391, 0.01151772, 0.01092881, 0.01092881, 0.01151772, 
    0.01180391, 0.001642336, 0,
  0, 0.01412936, 0.01151772, 0.006364421, 0.002450531, 0.002450531, 
    0.006364421, 0.01151772, 0.01412936, 0,
  0.002910513, 0.01096149, 0.01092881, 0.002450531, 0.00019574, 0.00019574, 
    0.002450531, 0.01092881, 0.01096149, 0.002910513,
  0.002910513, 0.01096149, 0.01092881, 0.002450531, 0.00019574, 0.00019574, 
    0.002450531, 0.01092881, 0.01096149, 0.002910513,
  0, 0.01412936, 0.01151772, 0.006364421, 0.002450531, 0.002450531, 
    0.006364421, 0.01151772, 0.01412936, 0,
  0, 0.001642336, 0.01180391, 0.01151772, 0.01092881, 0.01092881, 0.01151772, 
    0.01180391, 0.001642336, 0,
  0, 0, 0.001642336, 0.01412936, 0.01096149, 0.01096149, 0.01412936, 
    0.001642336, 0, 0,
  0, 0, 0, 0, 0.002910513, 0.002910513, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002905976, 0.002905976, 0, 0, 0, 0,
  0, 0, 0.00171827, 0.01403642, 0.01089066, 0.01089066, 0.01403642, 
    0.00171827, 0, 0,
  0, 0.00171827, 0.01170772, 0.01141188, 0.01082207, 0.01082207, 0.01141188, 
    0.01170772, 0.00171827, 0,
  0, 0.01403642, 0.01141188, 0.006238841, 0.002361601, 0.002361601, 
    0.006238841, 0.01141188, 0.01403642, 0,
  0.002905976, 0.01089066, 0.01082207, 0.002361601, 0.0001878417, 
    0.0001878417, 0.002361601, 0.01082207, 0.01089066, 0.002905976,
  0.002905976, 0.01089066, 0.01082207, 0.002361601, 0.0001878417, 
    0.0001878417, 0.002361601, 0.01082207, 0.01089066, 0.002905976,
  0, 0.01403642, 0.01141188, 0.006238841, 0.002361601, 0.002361601, 
    0.006238841, 0.01141188, 0.01403642, 0,
  0, 0.00171827, 0.01170772, 0.01141188, 0.01082207, 0.01082207, 0.01141188, 
    0.01170772, 0.00171827, 0,
  0, 0, 0.00171827, 0.01403642, 0.01089066, 0.01089066, 0.01403642, 
    0.00171827, 0, 0,
  0, 0, 0, 0, 0.002905976, 0.002905976, 0, 0, 0, 0,
  0, 0, 0, 0, 0.00281526, 0.00281526, 0, 0, 0, 0,
  0, 0, 0.00181455, 0.01361504, 0.01052553, 0.01052553, 0.01361504, 
    0.00181455, 0, 0,
  0, 0.00181455, 0.0113377, 0.01101774, 0.01039378, 0.01039378, 0.01101774, 
    0.0113377, 0.00181455, 0,
  0, 0.01361504, 0.01101774, 0.00589671, 0.002156245, 0.002156245, 
    0.00589671, 0.01101774, 0.01361504, 0,
  0.00281526, 0.01052553, 0.01039378, 0.002156245, 0.0001678793, 
    0.0001678793, 0.002156245, 0.01039378, 0.01052553, 0.00281526,
  0.00281526, 0.01052553, 0.01039378, 0.002156245, 0.0001678793, 
    0.0001678793, 0.002156245, 0.01039378, 0.01052553, 0.00281526,
  0, 0.01361504, 0.01101774, 0.00589671, 0.002156245, 0.002156245, 
    0.00589671, 0.01101774, 0.01361504, 0,
  0, 0.00181455, 0.0113377, 0.01101774, 0.01039378, 0.01039378, 0.01101774, 
    0.0113377, 0.00181455, 0,
  0, 0, 0.00181455, 0.01361504, 0.01052553, 0.01052553, 0.01361504, 
    0.00181455, 0, 0,
  0, 0, 0, 0, 0.00281526, 0.00281526, 0, 0, 0, 0,
  0, 0, 0, 0, 0.00259699, 0.00259699, 0, 0, 0, 0,
  0, 0, 0.001798689, 0.01259054, 0.009699423, 0.009699423, 0.01259054, 
    0.001798689, 0, 0,
  0, 0.001798689, 0.01049099, 0.01016702, 0.009561722, 0.009561722, 
    0.01016702, 0.01049099, 0.001798689, 0,
  0, 0.01259054, 0.01016702, 0.005365333, 0.00189847, 0.00189847, 
    0.005365333, 0.01016702, 0.01259054, 0,
  0.00259699, 0.009699423, 0.009561722, 0.00189847, 0.0001417474, 
    0.0001417474, 0.00189847, 0.009561722, 0.009699423, 0.00259699,
  0.00259699, 0.009699423, 0.009561722, 0.00189847, 0.0001417474, 
    0.0001417474, 0.00189847, 0.009561722, 0.009699423, 0.00259699,
  0, 0.01259054, 0.01016702, 0.005365333, 0.00189847, 0.00189847, 
    0.005365333, 0.01016702, 0.01259054, 0,
  0, 0.001798689, 0.01049099, 0.01016702, 0.009561722, 0.009561722, 
    0.01016702, 0.01049099, 0.001798689, 0,
  0, 0, 0.001798689, 0.01259054, 0.009699423, 0.009699423, 0.01259054, 
    0.001798689, 0, 0,
  0, 0, 0, 0, 0.00259699, 0.00259699, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002262004, 0.002262004, 0, 0, 0, 0,
  0, 0, 0.001653501, 0.01099986, 0.008444015, 0.008444015, 0.01099986, 
    0.001653501, 0, 0,
  0, 0.001653501, 0.009177292, 0.008872282, 0.008340399, 0.008340399, 
    0.008872282, 0.009177292, 0.001653501, 0,
  0, 0.01099986, 0.008872282, 0.004646091, 0.001606393, 0.001606393, 
    0.004646091, 0.008872282, 0.01099986, 0,
  0.002262004, 0.008444015, 0.008340399, 0.001606393, 0.0001149544, 
    0.0001149544, 0.001606393, 0.008340399, 0.008444015, 0.002262004,
  0.002262004, 0.008444015, 0.008340399, 0.001606393, 0.0001149544, 
    0.0001149544, 0.001606393, 0.008340399, 0.008444015, 0.002262004,
  0, 0.01099986, 0.008872282, 0.004646091, 0.001606393, 0.001606393, 
    0.004646091, 0.008872282, 0.01099986, 0,
  0, 0.001653501, 0.009177292, 0.008872282, 0.008340399, 0.008340399, 
    0.008872282, 0.009177292, 0.001653501, 0,
  0, 0, 0.001653501, 0.01099986, 0.008444015, 0.008444015, 0.01099986, 
    0.001653501, 0, 0,
  0, 0, 0, 0, 0.002262004, 0.002262004, 0, 0, 0, 0,
  0, 0, 0, 0, 0.001847901, 0.001847901, 0, 0, 0, 0,
  0, 0, 0.001407903, 0.009015079, 0.006896484, 0.006896484, 0.009015079, 
    0.001407903, 0, 0,
  0, 0.001407903, 0.007531525, 0.00726483, 0.006834279, 0.006834279, 
    0.00726483, 0.007531525, 0.001407903, 0,
  0, 0.009015079, 0.00726483, 0.003786854, 0.001289164, 0.001289164, 
    0.003786854, 0.00726483, 0.009015079, 0,
  0.001847901, 0.006896484, 0.006834279, 0.001289164, 8.961323e-05, 
    8.961323e-05, 0.001289164, 0.006834279, 0.006896484, 0.001847901,
  0.001847901, 0.006896484, 0.006834279, 0.001289164, 8.961323e-05, 
    8.961323e-05, 0.001289164, 0.006834279, 0.006896484, 0.001847901,
  0, 0.009015079, 0.00726483, 0.003786854, 0.001289164, 0.001289164, 
    0.003786854, 0.00726483, 0.009015079, 0,
  0, 0.001407903, 0.007531525, 0.00726483, 0.006834279, 0.006834279, 
    0.00726483, 0.007531525, 0.001407903, 0,
  0, 0, 0.001407903, 0.009015079, 0.006896484, 0.006896484, 0.009015079, 
    0.001407903, 0, 0,
  0, 0, 0, 0, 0.001847901, 0.001847901, 0, 0, 0, 0,
  0, 0, 0, 0, 0.001391239, 0.001391239, 0, 0, 0, 0,
  0, 0, 0.001095232, 0.00680995, 0.005191649, 0.005191649, 0.00680995, 
    0.001095232, 0, 0,
  0, 0.001095232, 0.00569629, 0.00548266, 0.005163534, 0.005163534, 
    0.00548266, 0.00569629, 0.001095232, 0,
  0, 0.00680995, 0.00548266, 0.002848994, 0.00095936, 0.00095936, 
    0.002848994, 0.00548266, 0.00680995, 0,
  0.001391239, 0.005191649, 0.005163534, 0.00095936, 6.562942e-05, 
    6.562942e-05, 0.00095936, 0.005163534, 0.005191649, 0.001391239,
  0.001391239, 0.005191649, 0.005163534, 0.00095936, 6.562942e-05, 
    6.562942e-05, 0.00095936, 0.005163534, 0.005191649, 0.001391239,
  0, 0.00680995, 0.00548266, 0.002848994, 0.00095936, 0.00095936, 
    0.002848994, 0.00548266, 0.00680995, 0,
  0, 0.001095232, 0.00569629, 0.00548266, 0.005163534, 0.005163534, 
    0.00548266, 0.00569629, 0.001095232, 0,
  0, 0, 0.001095232, 0.00680995, 0.005191649, 0.005191649, 0.00680995, 
    0.001095232, 0, 0,
  0, 0, 0, 0, 0.001391239, 0.001391239, 0, 0, 0, 0,
  0, 0, 0, 0, 0.000919933, 0.000919933, 0, 0, 0, 0,
  0, 0, 0.0007437959, 0.004519962, 0.003432815, 0.003432815, 0.004519962, 
    0.0007437959, 0, 0,
  0, 0.0007437959, 0.003784651, 0.003634558, 0.003427152, 0.003427152, 
    0.003634558, 0.003784651, 0.0007437959, 0,
  0, 0.004519962, 0.003634558, 0.001883997, 0.0006292354, 0.0006292354, 
    0.001883997, 0.003634558, 0.004519962, 0,
  0.000919933, 0.003432815, 0.003427152, 0.0006292354, 4.273657e-05, 
    4.273657e-05, 0.0006292354, 0.003427152, 0.003432815, 0.000919933,
  0.000919933, 0.003432815, 0.003427152, 0.0006292354, 4.273657e-05, 
    4.273657e-05, 0.0006292354, 0.003427152, 0.003432815, 0.000919933,
  0, 0.004519962, 0.003634558, 0.001883997, 0.0006292354, 0.0006292354, 
    0.001883997, 0.003634558, 0.004519962, 0,
  0, 0.0007437959, 0.003784651, 0.003634558, 0.003427152, 0.003427152, 
    0.003634558, 0.003784651, 0.0007437959, 0,
  0, 0, 0.0007437959, 0.004519962, 0.003432815, 0.003432815, 0.004519962, 
    0.0007437959, 0, 0,
  0, 0, 0, 0, 0.000919933, 0.000919933, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0004528118, 0.0004528118, 0, 0, 0, 0,
  0, 0, 0.0003748017, 0.002235653, 0.001689769, 0.001689769, 0.002235653, 
    0.0003748017, 0, 0,
  0, 0.0003748017, 0.001873085, 0.001794807, 0.001694755, 0.001694755, 
    0.001794807, 0.001873085, 0.0003748017, 0,
  0, 0.002235653, 0.001794807, 0.0009283751, 0.0003079593, 0.0003079593, 
    0.0009283751, 0.001794807, 0.002235653, 0,
  0.0004528118, 0.001689769, 0.001694755, 0.0003079593, 2.089243e-05, 
    2.089243e-05, 0.0003079593, 0.001694755, 0.001689769, 0.0004528118,
  0.0004528118, 0.001689769, 0.001694755, 0.0003079593, 2.089243e-05, 
    2.089243e-05, 0.0003079593, 0.001694755, 0.001689769, 0.0004528118,
  0, 0.002235653, 0.001794807, 0.0009283751, 0.0003079593, 0.0003079593, 
    0.0009283751, 0.001794807, 0.002235653, 0,
  0, 0.0003748017, 0.001873085, 0.001794807, 0.001694755, 0.001694755, 
    0.001794807, 0.001873085, 0.0003748017, 0,
  0, 0, 0.0003748017, 0.002235653, 0.001689769, 0.001689769, 0.002235653, 
    0.0003748017, 0, 0,
  0, 0, 0, 0, 0.0004528118, 0.0004528118, 0, 0, 0, 0,
  0, 0, 0, 0, 8.226774e-09, 8.226774e-09, 0, 0, 0, 0,
  0, 0, 1.730358e-08, 3.455538e-08, 3.655215e-08, 3.655215e-08, 3.455538e-08, 
    1.730358e-08, 0, 0,
  0, 1.730358e-08, 3.312687e-08, 2.959055e-08, 2.644049e-08, 2.644049e-08, 
    2.959055e-08, 3.312687e-08, 1.730358e-08, 0,
  0, 3.455538e-08, 2.959055e-08, 2.181365e-08, 1.611779e-08, 1.611779e-08, 
    2.181365e-08, 2.959055e-08, 3.455538e-08, 0,
  8.226774e-09, 3.655215e-08, 2.644049e-08, 1.611779e-08, 8.111424e-09, 
    8.111424e-09, 1.611779e-08, 2.644049e-08, 3.655215e-08, 8.226774e-09,
  8.226774e-09, 3.655215e-08, 2.644049e-08, 1.611779e-08, 8.111424e-09, 
    8.111424e-09, 1.611779e-08, 2.644049e-08, 3.655215e-08, 8.226774e-09,
  0, 3.455538e-08, 2.959055e-08, 2.181365e-08, 1.611779e-08, 1.611779e-08, 
    2.181365e-08, 2.959055e-08, 3.455538e-08, 0,
  0, 1.730358e-08, 3.312687e-08, 2.959055e-08, 2.644049e-08, 2.644049e-08, 
    2.959055e-08, 3.312687e-08, 1.730358e-08, 0,
  0, 0, 1.730358e-08, 3.455538e-08, 3.655215e-08, 3.655215e-08, 3.455538e-08, 
    1.730358e-08, 0, 0,
  0, 0, 0, 0, 8.226774e-09, 8.226774e-09, 0, 0, 0, 0,
  0, 0, 0, 0.0005935252, 0.0009224602, 0.0009224602, 0.0005935252, 0, 0, 0,
  0, 0, 0.0007205742, 0.002213747, 0.003449048, 0.003449048, 0.002213747, 
    0.0007205742, 0, 0,
  0, 0.0007205742, 0.0117114, 0.01093531, 0.009897564, 0.009897564, 
    0.01093531, 0.0117114, 0.0007205742, 0,
  0.0005935252, 0.002213747, 0.01093531, 0.006520234, 0.002520499, 
    0.002520499, 0.006520234, 0.01093531, 0.002213747, 0.0005935252,
  0.0009224602, 0.003449048, 0.009897564, 0.002520499, 0.0001945704, 
    0.0001945704, 0.002520499, 0.009897564, 0.003449048, 0.0009224602,
  0.0009224602, 0.003449048, 0.009897564, 0.002520499, 0.0001945704, 
    0.0001945704, 0.002520499, 0.009897564, 0.003449048, 0.0009224602,
  0.0005935252, 0.002213747, 0.01093531, 0.006520234, 0.002520499, 
    0.002520499, 0.006520234, 0.01093531, 0.002213747, 0.0005935252,
  0, 0.0007205742, 0.0117114, 0.01093531, 0.009897564, 0.009897564, 
    0.01093531, 0.0117114, 0.0007205742, 0,
  0, 0, 0.0007205742, 0.002213747, 0.003449048, 0.003449048, 0.002213747, 
    0.0007205742, 0, 0,
  0, 0, 0, 0.0005935252, 0.0009224602, 0.0009224602, 0.0005935252, 0, 0, 0,
  0, 0, 0, 0.00058077, 0.0009109076, 0.0009109076, 0.00058077, 0, 0, 0,
  0, 0, 0.0006429126, 0.002166014, 0.003401653, 0.003401653, 0.002166014, 
    0.0006429126, 0, 0,
  0, 0.0006429126, 0.01161182, 0.01081461, 0.009763596, 0.009763596, 
    0.01081461, 0.01161182, 0.0006429126, 0,
  0.00058077, 0.002166014, 0.01081461, 0.006410616, 0.002439159, 0.002439159, 
    0.006410616, 0.01081461, 0.002166014, 0.00058077,
  0.0009109076, 0.003401653, 0.009763596, 0.002439159, 0.0001830509, 
    0.0001830509, 0.002439159, 0.009763596, 0.003401653, 0.0009109076,
  0.0009109076, 0.003401653, 0.009763596, 0.002439159, 0.0001830509, 
    0.0001830509, 0.002439159, 0.009763596, 0.003401653, 0.0009109076,
  0.00058077, 0.002166014, 0.01081461, 0.006410616, 0.002439159, 0.002439159, 
    0.006410616, 0.01081461, 0.002166014, 0.00058077,
  0, 0.0006429126, 0.01161182, 0.01081461, 0.009763596, 0.009763596, 
    0.01081461, 0.01161182, 0.0006429126, 0,
  0, 0, 0.0006429126, 0.002166014, 0.003401653, 0.003401653, 0.002166014, 
    0.0006429126, 0, 0,
  0, 0, 0, 0.00058077, 0.0009109076, 0.0009109076, 0.00058077, 0, 0, 0,
  0, 0, 0, 0.0005484293, 0.0008751827, 0.0008751827, 0.0005484293, 0, 0, 0,
  0, 0, 0.0005070598, 0.002045693, 0.003266094, 0.003266094, 0.002045693, 
    0.0005070598, 0, 0,
  0, 0.0005070598, 0.01123223, 0.01043807, 0.009377853, 0.009377853, 
    0.01043807, 0.01123223, 0.0005070598, 0,
  0.0005484293, 0.002045693, 0.01043807, 0.006076507, 0.00223599, 0.00223599, 
    0.006076507, 0.01043807, 0.002045693, 0.0005484293,
  0.0008751827, 0.003266094, 0.009377853, 0.00223599, 0.0001604238, 
    0.0001604238, 0.00223599, 0.009377853, 0.003266094, 0.0008751827,
  0.0008751827, 0.003266094, 0.009377853, 0.00223599, 0.0001604238, 
    0.0001604238, 0.00223599, 0.009377853, 0.003266094, 0.0008751827,
  0.0005484293, 0.002045693, 0.01043807, 0.006076507, 0.00223599, 0.00223599, 
    0.006076507, 0.01043807, 0.002045693, 0.0005484293,
  0, 0.0005070598, 0.01123223, 0.01043807, 0.009377853, 0.009377853, 
    0.01043807, 0.01123223, 0.0005070598, 0,
  0, 0, 0.0005070598, 0.002045693, 0.003266094, 0.003266094, 0.002045693, 
    0.0005070598, 0, 0,
  0, 0, 0, 0.0005484293, 0.0008751827, 0.0008751827, 0.0005484293, 0, 0, 0,
  0, 0, 0, 0.0004957198, 0.0008012442, 0.0008012442, 0.0004957198, 0, 0, 0,
  0, 0, 0.000381839, 0.001849095, 0.0029894, 0.0029894, 0.001849095, 
    0.000381839, 0, 0,
  0, 0.000381839, 0.0103764, 0.009655268, 0.008655817, 0.008655817, 
    0.009655268, 0.0103764, 0.000381839, 0,
  0.0004957198, 0.001849095, 0.009655268, 0.00553204, 0.001972653, 
    0.001972653, 0.00553204, 0.009655268, 0.001849095, 0.0004957198,
  0.0008012442, 0.0029894, 0.008655817, 0.001972653, 0.0001335811, 
    0.0001335811, 0.001972653, 0.008655817, 0.0029894, 0.0008012442,
  0.0008012442, 0.0029894, 0.008655817, 0.001972653, 0.0001335811, 
    0.0001335811, 0.001972653, 0.008655817, 0.0029894, 0.0008012442,
  0.0004957198, 0.001849095, 0.009655268, 0.00553204, 0.001972653, 
    0.001972653, 0.00553204, 0.009655268, 0.001849095, 0.0004957198,
  0, 0.000381839, 0.0103764, 0.009655268, 0.008655817, 0.008655817, 
    0.009655268, 0.0103764, 0.000381839, 0,
  0, 0, 0.000381839, 0.001849095, 0.0029894, 0.0029894, 0.001849095, 
    0.000381839, 0, 0,
  0, 0, 0, 0.0004957198, 0.0008012442, 0.0008012442, 0.0004957198, 0, 0, 0,
  0, 0, 0, 0.0004250235, 0.0006929337, 0.0006929337, 0.0004250235, 0, 0, 0,
  0, 0, 0.000278449, 0.001585442, 0.002585121, 0.002585121, 0.001585442, 
    0.000278449, 0, 0,
  0, 0.000278449, 0.00906265, 0.008453338, 0.007580093, 0.007580093, 
    0.008453338, 0.00906265, 0.000278449, 0,
  0.0004250235, 0.001585442, 0.008453338, 0.004787584, 0.001670079, 
    0.001670079, 0.004787584, 0.008453338, 0.001585442, 0.0004250235,
  0.0006929337, 0.002585121, 0.007580093, 0.001670079, 0.000107436, 
    0.000107436, 0.001670079, 0.007580093, 0.002585121, 0.0006929337,
  0.0006929337, 0.002585121, 0.007580093, 0.001670079, 0.000107436, 
    0.000107436, 0.001670079, 0.007580093, 0.002585121, 0.0006929337,
  0.0004250235, 0.001585442, 0.008453338, 0.004787584, 0.001670079, 
    0.001670079, 0.004787584, 0.008453338, 0.001585442, 0.0004250235,
  0, 0.000278449, 0.00906265, 0.008453338, 0.007580093, 0.007580093, 
    0.008453338, 0.00906265, 0.000278449, 0,
  0, 0, 0.000278449, 0.001585442, 0.002585121, 0.002585121, 0.001585442, 
    0.000278449, 0, 0,
  0, 0, 0, 0.0004250235, 0.0006929337, 0.0006929337, 0.0004250235, 0, 0, 0,
  0, 0, 0, 0.0003429074, 0.0005625431, 0.0005625431, 0.0003429074, 0, 0, 0,
  0, 0, 0.000195564, 0.001279208, 0.002098703, 0.002098703, 0.001279208, 
    0.000195564, 0, 0,
  0, 0.000195564, 0.007427904, 0.006944943, 0.006234465, 0.006234465, 
    0.006944943, 0.007427904, 0.000195564, 0,
  0.0003429074, 0.001279208, 0.006944943, 0.003898633, 0.001340065, 
    0.001340065, 0.003898633, 0.006944943, 0.001279208, 0.0003429074,
  0.0005625431, 0.002098703, 0.006234465, 0.001340065, 8.343284e-05, 
    8.343284e-05, 0.001340065, 0.006234465, 0.002098703, 0.0005625431,
  0.0005625431, 0.002098703, 0.006234465, 0.001340065, 8.343284e-05, 
    8.343284e-05, 0.001340065, 0.006234465, 0.002098703, 0.0005625431,
  0.0003429074, 0.001279208, 0.006944943, 0.003898633, 0.001340065, 
    0.001340065, 0.003898633, 0.006944943, 0.001279208, 0.0003429074,
  0, 0.000195564, 0.007427904, 0.006944943, 0.006234465, 0.006234465, 
    0.006944943, 0.007427904, 0.000195564, 0,
  0, 0, 0.000195564, 0.001279208, 0.002098703, 0.002098703, 0.001279208, 
    0.000195564, 0, 0,
  0, 0, 0, 0.0003429074, 0.0005625431, 0.0005625431, 0.0003429074, 0, 0, 0,
  0, 0, 0, 0.0002556448, 0.0004212726, 0.0004212726, 0.0002556448, 0, 0, 0,
  0, 0, 0.0001303855, 0.0009537524, 0.001571744, 0.001571744, 0.0009537524, 
    0.0001303855, 0, 0,
  0, 0.0001303855, 0.005613131, 0.005258332, 0.004726373, 0.004726373, 
    0.005258332, 0.005613131, 0.0001303855, 0,
  0.0002556448, 0.0009537524, 0.005258332, 0.002930569, 0.000996945, 
    0.000996945, 0.002930569, 0.005258332, 0.0009537524, 0.0002556448,
  0.0004212726, 0.001571744, 0.004726373, 0.000996945, 6.103645e-05, 
    6.103645e-05, 0.000996945, 0.004726373, 0.001571744, 0.0004212726,
  0.0004212726, 0.001571744, 0.004726373, 0.000996945, 6.103645e-05, 
    6.103645e-05, 0.000996945, 0.004726373, 0.001571744, 0.0004212726,
  0.0002556448, 0.0009537524, 0.005258332, 0.002930569, 0.000996945, 
    0.000996945, 0.002930569, 0.005258332, 0.0009537524, 0.0002556448,
  0, 0.0001303855, 0.005613131, 0.005258332, 0.004726373, 0.004726373, 
    0.005258332, 0.005613131, 0.0001303855, 0,
  0, 0, 0.0001303855, 0.0009537524, 0.001571744, 0.001571744, 0.0009537524, 
    0.0001303855, 0, 0,
  0, 0, 0, 0.0002556448, 0.0004212726, 0.0004212726, 0.0002556448, 0, 0, 0,
  0, 0, 0, 0.0001677808, 0.0002773091, 0.0002773091, 0.0001677808, 0, 0, 0,
  0, 0, 7.884818e-05, 0.0006260082, 0.001034704, 0.001034704, 0.0006260082, 
    7.884818e-05, 0, 0,
  0, 7.884818e-05, 0.003728302, 0.003497615, 0.003147299, 0.003147299, 
    0.003497615, 0.003728302, 7.884818e-05, 0,
  0.0001677808, 0.0006260082, 0.003497615, 0.001936881, 0.0006538513, 
    0.0006538513, 0.001936881, 0.003497615, 0.0006260082, 0.0001677808,
  0.0002773091, 0.001034704, 0.003147299, 0.0006538513, 3.976773e-05, 
    3.976773e-05, 0.0006538513, 0.003147299, 0.001034704, 0.0002773091,
  0.0002773091, 0.001034704, 0.003147299, 0.0006538513, 3.976773e-05, 
    3.976773e-05, 0.0006538513, 0.003147299, 0.001034704, 0.0002773091,
  0.0001677808, 0.0006260082, 0.003497615, 0.001936881, 0.0006538513, 
    0.0006538513, 0.001936881, 0.003497615, 0.0006260082, 0.0001677808,
  0, 7.884818e-05, 0.003728302, 0.003497615, 0.003147299, 0.003147299, 
    0.003497615, 0.003728302, 7.884818e-05, 0,
  0, 0, 7.884818e-05, 0.0006260082, 0.001034704, 0.001034704, 0.0006260082, 
    7.884818e-05, 0, 0,
  0, 0, 0, 0.0001677808, 0.0002773091, 0.0002773091, 0.0001677808, 0, 0, 0,
  0, 0, 0, 8.210483e-05, 0.0001359555, 0.0001359555, 8.210483e-05, 0, 0, 0,
  0, 0, 3.6514e-05, 0.0003063745, 0.0005073319, 0.0005073319, 0.0003063745, 
    3.6514e-05, 0, 0,
  0, 3.6514e-05, 0.001845718, 0.001734024, 0.001562124, 0.001562124, 
    0.001734024, 0.001845718, 3.6514e-05, 0,
  8.210483e-05, 0.0003063745, 0.001734024, 0.0009548268, 0.000320278, 
    0.000320278, 0.0009548268, 0.001734024, 0.0003063745, 8.210483e-05,
  0.0001359555, 0.0005073319, 0.001562124, 0.000320278, 1.947795e-05, 
    1.947795e-05, 0.000320278, 0.001562124, 0.0005073319, 0.0001359555,
  0.0001359555, 0.0005073319, 0.001562124, 0.000320278, 1.947795e-05, 
    1.947795e-05, 0.000320278, 0.001562124, 0.0005073319, 0.0001359555,
  8.210483e-05, 0.0003063745, 0.001734024, 0.0009548268, 0.000320278, 
    0.000320278, 0.0009548268, 0.001734024, 0.0003063745, 8.210483e-05,
  0, 3.6514e-05, 0.001845718, 0.001734024, 0.001562124, 0.001562124, 
    0.001734024, 0.001845718, 3.6514e-05, 0,
  0, 0, 3.6514e-05, 0.0003063745, 0.0005073319, 0.0005073319, 0.0003063745, 
    3.6514e-05, 0, 0,
  0, 0, 0, 8.210483e-05, 0.0001359555, 0.0001359555, 8.210483e-05, 0, 0, 0,
  0, 0, 0, 5.83815e-09, 7.008377e-09, 7.008377e-09, 5.83815e-09, 0, 0, 0,
  0, 0, 1.751749e-08, 2.412821e-08, 2.865664e-08, 2.865664e-08, 2.412821e-08, 
    1.751749e-08, 0, 0,
  0, 1.751749e-08, 3.31963e-08, 2.920203e-08, 2.597933e-08, 2.597933e-08, 
    2.920203e-08, 3.31963e-08, 1.751749e-08, 0,
  5.83815e-09, 2.412821e-08, 2.920203e-08, 2.183868e-08, 1.61319e-08, 
    1.61319e-08, 2.183868e-08, 2.920203e-08, 2.412821e-08, 5.83815e-09,
  7.008377e-09, 2.865664e-08, 2.597933e-08, 1.61319e-08, 8.202348e-09, 
    8.202348e-09, 1.61319e-08, 2.597933e-08, 2.865664e-08, 7.008377e-09,
  7.008377e-09, 2.865664e-08, 2.597933e-08, 1.61319e-08, 8.202348e-09, 
    8.202348e-09, 1.61319e-08, 2.597933e-08, 2.865664e-08, 7.008377e-09,
  5.83815e-09, 2.412821e-08, 2.920203e-08, 2.183868e-08, 1.61319e-08, 
    1.61319e-08, 2.183868e-08, 2.920203e-08, 2.412821e-08, 5.83815e-09,
  0, 1.751749e-08, 3.31963e-08, 2.920203e-08, 2.597933e-08, 2.597933e-08, 
    2.920203e-08, 3.31963e-08, 1.751749e-08, 0,
  0, 0, 1.751749e-08, 2.412821e-08, 2.865664e-08, 2.865664e-08, 2.412821e-08, 
    1.751749e-08, 0, 0,
  0, 0, 0, 5.83815e-09, 7.008377e-09, 7.008377e-09, 5.83815e-09, 0, 0, 0,
  0, 0, 0, 0.0005984311, 0.0009270075, 0.0009270075, 0.0005984311, 0, 0, 0,
  0, 0, 0.0007392654, 0.002232191, 0.0034662, 0.0034662, 0.002232191, 
    0.0007392654, 0, 0,
  0, 0.0007392654, 0.01172141, 0.01089894, 0.009836782, 0.009836782, 
    0.01089894, 0.01172141, 0.0007392654, 0,
  0.0005984311, 0.002232191, 0.01089894, 0.006497891, 0.002526133, 
    0.002526133, 0.006497891, 0.01089894, 0.002232191, 0.0005984311,
  0.0009270075, 0.0034662, 0.009836782, 0.002526133, 0.0001981906, 
    0.0001981906, 0.002526133, 0.009836782, 0.0034662, 0.0009270075,
  0.0009270075, 0.0034662, 0.009836782, 0.002526133, 0.0001981906, 
    0.0001981906, 0.002526133, 0.009836782, 0.0034662, 0.0009270075,
  0.0005984311, 0.002232191, 0.01089894, 0.006497891, 0.002526133, 
    0.002526133, 0.006497891, 0.01089894, 0.002232191, 0.0005984311,
  0, 0.0007392654, 0.01172141, 0.01089894, 0.009836782, 0.009836782, 
    0.01089894, 0.01172141, 0.0007392654, 0,
  0, 0, 0.0007392654, 0.002232191, 0.0034662, 0.0034662, 0.002232191, 
    0.0007392654, 0, 0,
  0, 0, 0, 0.0005984311, 0.0009270075, 0.0009270075, 0.0005984311, 0, 0, 0,
  0, 0, 0, 0.0005856783, 0.0009154733, 0.0009154733, 0.0005856783, 0, 0, 0,
  0, 0, 0.0006615929, 0.002184406, 0.003418792, 0.003418792, 0.002184406, 
    0.0006615929, 0, 0,
  0, 0.0006615929, 0.01162179, 0.01077886, 0.00970428, 0.00970428, 
    0.01077886, 0.01162179, 0.0006615929, 0,
  0.0005856783, 0.002184406, 0.01077886, 0.006388575, 0.002444883, 
    0.002444883, 0.006388575, 0.01077886, 0.002184406, 0.0005856783,
  0.0009154733, 0.003418792, 0.00970428, 0.002444883, 0.000186501, 
    0.000186501, 0.002444883, 0.00970428, 0.003418792, 0.0009154733,
  0.0009154733, 0.003418792, 0.00970428, 0.002444883, 0.000186501, 
    0.000186501, 0.002444883, 0.00970428, 0.003418792, 0.0009154733,
  0.0005856783, 0.002184406, 0.01077886, 0.006388575, 0.002444883, 
    0.002444883, 0.006388575, 0.01077886, 0.002184406, 0.0005856783,
  0, 0.0006615929, 0.01162179, 0.01077886, 0.00970428, 0.00970428, 
    0.01077886, 0.01162179, 0.0006615929, 0,
  0, 0, 0.0006615929, 0.002184406, 0.003418792, 0.003418792, 0.002184406, 
    0.0006615929, 0, 0,
  0, 0, 0, 0.0005856783, 0.0009154733, 0.0009154733, 0.0005856783, 0, 0, 0,
  0, 0, 0, 0.0005532826, 0.0008796834, 0.0008796834, 0.0005532826, 0, 0, 0,
  0, 0, 0.0005249733, 0.002063841, 0.00328294, 0.00328294, 0.002063841, 
    0.0005249733, 0, 0,
  0, 0.0005249733, 0.01124249, 0.010404, 0.009321776, 0.009321776, 0.010404, 
    0.01124249, 0.0005249733, 0,
  0.0005532826, 0.002063841, 0.010404, 0.006055712, 0.002242041, 0.002242041, 
    0.006055712, 0.010404, 0.002063841, 0.0005532826,
  0.0008796834, 0.00328294, 0.009321776, 0.002242041, 0.0001634534, 
    0.0001634534, 0.002242041, 0.009321776, 0.00328294, 0.0008796834,
  0.0008796834, 0.00328294, 0.009321776, 0.002242041, 0.0001634534, 
    0.0001634534, 0.002242041, 0.009321776, 0.00328294, 0.0008796834,
  0.0005532826, 0.002063841, 0.010404, 0.006055712, 0.002242041, 0.002242041, 
    0.006055712, 0.010404, 0.002063841, 0.0005532826,
  0, 0.0005249733, 0.01124249, 0.010404, 0.009321776, 0.009321776, 0.010404, 
    0.01124249, 0.0005249733, 0,
  0, 0, 0.0005249733, 0.002063841, 0.00328294, 0.00328294, 0.002063841, 
    0.0005249733, 0, 0,
  0, 0, 0, 0.0005532826, 0.0008796834, 0.0008796834, 0.0005532826, 0, 0, 0,
  0, 0, 0, 0.000500294, 0.0008054702, 0.0008054702, 0.000500294, 0, 0, 0,
  0, 0, 0.0003979405, 0.001866183, 0.003005198, 0.003005198, 0.001866183, 
    0.0003979405, 0, 0,
  0, 0.0003979405, 0.01038728, 0.009624528, 0.008604906, 0.008604906, 
    0.009624528, 0.01038728, 0.0003979405, 0,
  0.000500294, 0.001866183, 0.009624528, 0.005513341, 0.001978825, 
    0.001978825, 0.005513341, 0.009624528, 0.001866183, 0.000500294,
  0.0008054702, 0.003005198, 0.008604906, 0.001978825, 0.0001361242, 
    0.0001361242, 0.001978825, 0.008604906, 0.003005198, 0.0008054702,
  0.0008054702, 0.003005198, 0.008604906, 0.001978825, 0.0001361242, 
    0.0001361242, 0.001978825, 0.008604906, 0.003005198, 0.0008054702,
  0.000500294, 0.001866183, 0.009624528, 0.005513341, 0.001978825, 
    0.001978825, 0.005513341, 0.009624528, 0.001866183, 0.000500294,
  0, 0.0003979405, 0.01038728, 0.009624528, 0.008604906, 0.008604906, 
    0.009624528, 0.01038728, 0.0003979405, 0,
  0, 0, 0.0003979405, 0.001866183, 0.003005198, 0.003005198, 0.001866183, 
    0.0003979405, 0, 0,
  0, 0, 0, 0.000500294, 0.0008054702, 0.0008054702, 0.000500294, 0, 0, 0,
  0, 0, 0, 0.0004291001, 0.0006966924, 0.0006966924, 0.0004291001, 0, 0, 0,
  0, 0, 0.0002919014, 0.001600663, 0.002599162, 0.002599162, 0.001600663, 
    0.0002919014, 0, 0,
  0, 0.0002919014, 0.009074253, 0.008427681, 0.007536518, 0.007536518, 
    0.008427681, 0.009074253, 0.0002919014, 0,
  0.0004291001, 0.001600663, 0.008427681, 0.004771727, 0.001675924, 
    0.001675924, 0.004771727, 0.008427681, 0.001600663, 0.0004291001,
  0.0006966924, 0.002599162, 0.007536518, 0.001675924, 0.0001095178, 
    0.0001095178, 0.001675924, 0.007536518, 0.002599162, 0.0006966924,
  0.0006966924, 0.002599162, 0.007536518, 0.001675924, 0.0001095178, 
    0.0001095178, 0.001675924, 0.007536518, 0.002599162, 0.0006966924,
  0.0004291001, 0.001600663, 0.008427681, 0.004771727, 0.001675924, 
    0.001675924, 0.004771727, 0.008427681, 0.001600663, 0.0004291001,
  0, 0.0002919014, 0.009074253, 0.008427681, 0.007536518, 0.007536518, 
    0.008427681, 0.009074253, 0.0002919014, 0,
  0, 0, 0.0002919014, 0.001600663, 0.002599162, 0.002599162, 0.001600663, 
    0.0002919014, 0, 0,
  0, 0, 0, 0.0004291001, 0.0006966924, 0.0006966924, 0.0004291001, 0, 0, 0,
  0, 0, 0, 0.000346336, 0.0005656932, 0.0005656932, 0.000346336, 0, 0, 0,
  0, 0, 0.0002059765, 0.001292006, 0.002110465, 0.002110465, 0.001292006, 
    0.0002059765, 0, 0,
  0, 0.0002059765, 0.007440123, 0.006925647, 0.006199959, 0.006199959, 
    0.006925647, 0.007440123, 0.0002059765, 0,
  0.000346336, 0.001292006, 0.006925647, 0.003886177, 0.001345212, 
    0.001345212, 0.003886177, 0.006925647, 0.001292006, 0.000346336,
  0.0005656932, 0.002110465, 0.006199959, 0.001345212, 8.508114e-05, 
    8.508114e-05, 0.001345212, 0.006199959, 0.002110465, 0.0005656932,
  0.0005656932, 0.002110465, 0.006199959, 0.001345212, 8.508114e-05, 
    8.508114e-05, 0.001345212, 0.006199959, 0.002110465, 0.0005656932,
  0.000346336, 0.001292006, 0.006925647, 0.003886177, 0.001345212, 
    0.001345212, 0.003886177, 0.006925647, 0.001292006, 0.000346336,
  0, 0.0002059765, 0.007440123, 0.006925647, 0.006199959, 0.006199959, 
    0.006925647, 0.007440123, 0.0002059765, 0,
  0, 0, 0.0002059765, 0.001292006, 0.002110465, 0.002110465, 0.001292006, 
    0.0002059765, 0, 0,
  0, 0, 0, 0.000346336, 0.0005656932, 0.0005656932, 0.000346336, 0, 0, 0,
  0, 0, 0, 0.0002583319, 0.0004237273, 0.0004237273, 0.0002583319, 0, 0, 0,
  0, 0, 0.0001377579, 0.0009637799, 0.001580907, 0.001580907, 0.0009637799, 
    0.0001377579, 0, 0,
  0, 0.0001377579, 0.005625602, 0.005246054, 0.004701991, 0.004701991, 
    0.005246054, 0.005625602, 0.0001377579, 0,
  0.0002583319, 0.0009637799, 0.005246054, 0.002921861, 0.001001161, 
    0.001001161, 0.002921861, 0.005246054, 0.0009637799, 0.0002583319,
  0.0004237273, 0.001580907, 0.004701991, 0.001001161, 6.227034e-05, 
    6.227034e-05, 0.001001161, 0.004701991, 0.001580907, 0.0004237273,
  0.0004237273, 0.001580907, 0.004701991, 0.001001161, 6.227034e-05, 
    6.227034e-05, 0.001001161, 0.004701991, 0.001580907, 0.0004237273,
  0.0002583319, 0.0009637799, 0.005246054, 0.002921861, 0.001001161, 
    0.001001161, 0.002921861, 0.005246054, 0.0009637799, 0.0002583319,
  0, 0.0001377579, 0.005625602, 0.005246054, 0.004701991, 0.004701991, 
    0.005246054, 0.005625602, 0.0001377579, 0,
  0, 0, 0.0001377579, 0.0009637799, 0.001580907, 0.001580907, 0.0009637799, 
    0.0001377579, 0, 0,
  0, 0, 0, 0.0002583319, 0.0004237273, 0.0004237273, 0.0002583319, 0, 0, 0,
  0, 0, 0, 0.000169655, 0.0002790212, 0.0002790212, 0.000169655, 0, 0, 0,
  0, 0, 8.338108e-05, 0.0006330012, 0.001041093, 0.001041093, 0.0006330012, 
    8.338108e-05, 0, 0,
  0, 8.338108e-05, 0.003739877, 0.003492221, 0.003133371, 0.003133371, 
    0.003492221, 0.003739877, 8.338108e-05, 0,
  0.000169655, 0.0006330012, 0.003492221, 0.001932136, 0.0006570021, 
    0.0006570021, 0.001932136, 0.003492221, 0.0006330012, 0.000169655,
  0.0002790212, 0.001041093, 0.003133371, 0.0006570021, 4.060302e-05, 
    4.060302e-05, 0.0006570021, 0.003133371, 0.001041093, 0.0002790212,
  0.0002790212, 0.001041093, 0.003133371, 0.0006570021, 4.060302e-05, 
    4.060302e-05, 0.0006570021, 0.003133371, 0.001041093, 0.0002790212,
  0.000169655, 0.0006330012, 0.003492221, 0.001932136, 0.0006570021, 
    0.0006570021, 0.001932136, 0.003492221, 0.0006330012, 0.000169655,
  0, 8.338108e-05, 0.003739877, 0.003492221, 0.003133371, 0.003133371, 
    0.003492221, 0.003739877, 8.338108e-05, 0,
  0, 0, 8.338108e-05, 0.0006330012, 0.001041093, 0.001041093, 0.0006330012, 
    8.338108e-05, 0, 0,
  0, 0, 0, 0.000169655, 0.0002790212, 0.0002790212, 0.000169655, 0, 0, 0,
  0, 0, 0, 8.307464e-05, 0.0001368674, 0.0001368674, 8.307464e-05, 0, 0, 0,
  0, 0, 3.846741e-05, 0.0003099931, 0.0005107349, 0.0005107349, 0.0003099931, 
    3.846741e-05, 0, 0,
  0, 3.846741e-05, 0.001853527, 0.001733682, 0.001557494, 0.001557494, 
    0.001733682, 0.001853527, 3.846741e-05, 0,
  8.307464e-05, 0.0003099931, 0.001733682, 0.0009538077, 0.0003222257, 
    0.0003222257, 0.0009538077, 0.001733682, 0.0003099931, 8.307464e-05,
  0.0001368674, 0.0005107349, 0.001557494, 0.0003222257, 1.991739e-05, 
    1.991739e-05, 0.0003222257, 0.001557494, 0.0005107349, 0.0001368674,
  0.0001368674, 0.0005107349, 0.001557494, 0.0003222257, 1.991739e-05, 
    1.991739e-05, 0.0003222257, 0.001557494, 0.0005107349, 0.0001368674,
  8.307464e-05, 0.0003099931, 0.001733682, 0.0009538077, 0.0003222257, 
    0.0003222257, 0.0009538077, 0.001733682, 0.0003099931, 8.307464e-05,
  0, 3.846741e-05, 0.001853527, 0.001733682, 0.001557494, 0.001557494, 
    0.001733682, 0.001853527, 3.846741e-05, 0,
  0, 0, 3.846741e-05, 0.0003099931, 0.0005107349, 0.0005107349, 0.0003099931, 
    3.846741e-05, 0, 0,
  0, 0, 0, 8.307464e-05, 0.0001368674, 0.0001368674, 8.307464e-05, 0, 0, 0,
  0, 0, 0, 5.84133e-09, 7.008931e-09, 7.008931e-09, 5.84133e-09, 0, 0, 0,
  0, 0, 1.754809e-08, 2.415812e-08, 2.868049e-08, 2.868049e-08, 2.415812e-08, 
    1.754809e-08, 0, 0,
  0, 1.754809e-08, 3.31868e-08, 2.915244e-08, 2.590853e-08, 2.590853e-08, 
    2.915244e-08, 3.31868e-08, 1.754809e-08, 0,
  5.84133e-09, 2.415812e-08, 2.915244e-08, 2.181345e-08, 1.61398e-08, 
    1.61398e-08, 2.181345e-08, 2.915244e-08, 2.415812e-08, 5.84133e-09,
  7.008931e-09, 2.868049e-08, 2.590853e-08, 1.61398e-08, 8.232286e-09, 
    8.232286e-09, 1.61398e-08, 2.590853e-08, 2.868049e-08, 7.008931e-09,
  7.008931e-09, 2.868049e-08, 2.590853e-08, 1.61398e-08, 8.232286e-09, 
    8.232286e-09, 1.61398e-08, 2.590853e-08, 2.868049e-08, 7.008931e-09,
  5.84133e-09, 2.415812e-08, 2.915244e-08, 2.181345e-08, 1.61398e-08, 
    1.61398e-08, 2.181345e-08, 2.915244e-08, 2.415812e-08, 5.84133e-09,
  0, 1.754809e-08, 3.31868e-08, 2.915244e-08, 2.590853e-08, 2.590853e-08, 
    2.915244e-08, 3.31868e-08, 1.754809e-08, 0,
  0, 0, 1.754809e-08, 2.415812e-08, 2.868049e-08, 2.868049e-08, 2.415812e-08, 
    1.754809e-08, 0, 0,
  0, 0, 0, 5.84133e-09, 7.008931e-09, 7.008931e-09, 5.84133e-09, 0, 0, 0,
  0, 0, 0, 0.0006027271, 0.0009310155, 0.0009310155, 0.0006027271, 0, 0, 0,
  0, 0, 0.0007588615, 0.002248328, 0.003481323, 0.003481323, 0.002248328, 
    0.0007588615, 0, 0,
  0, 0.0007588615, 0.01173086, 0.01086331, 0.009777134, 0.009777134, 
    0.01086331, 0.01173086, 0.0007588615, 0,
  0.0006027271, 0.002248328, 0.01086331, 0.006475622, 0.002531606, 
    0.002531606, 0.006475622, 0.01086331, 0.002248328, 0.0006027271,
  0.0009310155, 0.003481323, 0.009777134, 0.002531606, 0.0002018188, 
    0.0002018188, 0.002531606, 0.009777134, 0.003481323, 0.0009310155,
  0.0009310155, 0.003481323, 0.009777134, 0.002531606, 0.0002018188, 
    0.0002018188, 0.002531606, 0.009777134, 0.003481323, 0.0009310155,
  0.0006027271, 0.002248328, 0.01086331, 0.006475622, 0.002531606, 
    0.002531606, 0.006475622, 0.01086331, 0.002248328, 0.0006027271,
  0, 0.0007588615, 0.01173086, 0.01086331, 0.009777134, 0.009777134, 
    0.01086331, 0.01173086, 0.0007588615, 0,
  0, 0, 0.0007588615, 0.002248328, 0.003481323, 0.003481323, 0.002248328, 
    0.0007588615, 0, 0,
  0, 0, 0, 0.0006027271, 0.0009310155, 0.0009310155, 0.0006027271, 0, 0, 0,
  0, 0, 0, 0.0005899783, 0.0009195007, 0.0009195007, 0.0005899783, 0, 0, 0,
  0, 0, 0.000681197, 0.002200501, 0.00343391, 0.00343391, 0.002200501, 
    0.000681197, 0, 0,
  0, 0.000681197, 0.01163121, 0.01074382, 0.009646049, 0.009646049, 
    0.01074382, 0.01163121, 0.000681197, 0,
  0.0005899783, 0.002200501, 0.01074382, 0.006366613, 0.002450452, 
    0.002450452, 0.006366613, 0.01074382, 0.002200501, 0.0005899783,
  0.0009195007, 0.00343391, 0.009646049, 0.002450452, 0.0001899589, 
    0.0001899589, 0.002450452, 0.009646049, 0.00343391, 0.0009195007,
  0.0009195007, 0.00343391, 0.009646049, 0.002450452, 0.0001899589, 
    0.0001899589, 0.002450452, 0.009646049, 0.00343391, 0.0009195007,
  0.0005899783, 0.002200501, 0.01074382, 0.006366613, 0.002450452, 
    0.002450452, 0.006366613, 0.01074382, 0.002200501, 0.0005899783,
  0, 0.000681197, 0.01163121, 0.01074382, 0.009646049, 0.009646049, 
    0.01074382, 0.01163121, 0.000681197, 0,
  0, 0, 0.000681197, 0.002200501, 0.00343391, 0.00343391, 0.002200501, 
    0.000681197, 0, 0,
  0, 0, 0, 0.0005899783, 0.0009195007, 0.0009195007, 0.0005899783, 0, 0, 0,
  0, 0, 0, 0.0005575338, 0.0008836526, 0.0008836526, 0.0005575338, 0, 0, 0,
  0, 0, 0.0005438611, 0.002079721, 0.003297795, 0.003297795, 0.002079721, 
    0.0005438611, 0, 0,
  0, 0.0005438611, 0.01125222, 0.01037059, 0.009266708, 0.009266708, 
    0.01037059, 0.01125222, 0.0005438611, 0,
  0.0005575338, 0.002079721, 0.01037059, 0.006034989, 0.002247942, 
    0.002247942, 0.006034989, 0.01037059, 0.002079721, 0.0005575338,
  0.0008836526, 0.003297795, 0.009266708, 0.002247942, 0.0001664922, 
    0.0001664922, 0.002247942, 0.009266708, 0.003297795, 0.0008836526,
  0.0008836526, 0.003297795, 0.009266708, 0.002247942, 0.0001664922, 
    0.0001664922, 0.002247942, 0.009266708, 0.003297795, 0.0008836526,
  0.0005575338, 0.002079721, 0.01037059, 0.006034989, 0.002247942, 
    0.002247942, 0.006034989, 0.01037059, 0.002079721, 0.0005575338,
  0, 0.0005438611, 0.01125222, 0.01037059, 0.009266708, 0.009266708, 
    0.01037059, 0.01125222, 0.0005438611, 0,
  0, 0, 0.0005438611, 0.002079721, 0.003297795, 0.003297795, 0.002079721, 
    0.0005438611, 0, 0,
  0, 0, 0, 0.0005575338, 0.0008836526, 0.0008836526, 0.0005575338, 0, 0, 0,
  0, 0, 0, 0.0005042931, 0.0008091935, 0.0008091935, 0.0005042931, 0, 0, 0,
  0, 0, 0.0004150518, 0.001881107, 0.003019114, 0.003019114, 0.001881107, 
    0.0004150518, 0, 0,
  0, 0.0004150518, 0.01039764, 0.009594386, 0.008554914, 0.008554914, 
    0.009594386, 0.01039764, 0.0004150518, 0,
  0.0005042931, 0.001881107, 0.009594386, 0.005494698, 0.001984854, 
    0.001984854, 0.005494698, 0.009594386, 0.001881107, 0.0005042931,
  0.0008091935, 0.003019114, 0.008554914, 0.001984854, 0.0001386789, 
    0.0001386789, 0.001984854, 0.008554914, 0.003019114, 0.0008091935,
  0.0008091935, 0.003019114, 0.008554914, 0.001984854, 0.0001386789, 
    0.0001386789, 0.001984854, 0.008554914, 0.003019114, 0.0008091935,
  0.0005042931, 0.001881107, 0.009594386, 0.005494698, 0.001984854, 
    0.001984854, 0.005494698, 0.009594386, 0.001881107, 0.0005042931,
  0, 0.0004150518, 0.01039764, 0.009594386, 0.008554914, 0.008554914, 
    0.009594386, 0.01039764, 0.0004150518, 0,
  0, 0, 0.0004150518, 0.001881107, 0.003019114, 0.003019114, 0.001881107, 
    0.0004150518, 0, 0,
  0, 0, 0, 0.0005042931, 0.0008091935, 0.0008091935, 0.0005042931, 0, 0, 0,
  0, 0, 0, 0.0004326566, 0.0007000027, 0.0007000027, 0.0004326566, 0, 0, 0,
  0, 0, 0.0003063596, 0.00161393, 0.002611525, 0.002611525, 0.00161393, 
    0.0003063596, 0, 0,
  0, 0.0003063596, 0.00908535, 0.008402547, 0.00749374, 0.00749374, 
    0.008402547, 0.00908535, 0.0003063596, 0,
  0.0004326566, 0.00161393, 0.008402547, 0.00475591, 0.001681639, 
    0.001681639, 0.00475591, 0.008402547, 0.00161393, 0.0004326566,
  0.0007000027, 0.002611525, 0.00749374, 0.001681639, 0.000111612, 
    0.000111612, 0.001681639, 0.00749374, 0.002611525, 0.0007000027,
  0.0007000027, 0.002611525, 0.00749374, 0.001681639, 0.000111612, 
    0.000111612, 0.001681639, 0.00749374, 0.002611525, 0.0007000027,
  0.0004326566, 0.00161393, 0.008402547, 0.00475591, 0.001681639, 
    0.001681639, 0.00475591, 0.008402547, 0.00161393, 0.0004326566,
  0, 0.0003063596, 0.00908535, 0.008402547, 0.00749374, 0.00749374, 
    0.008402547, 0.00908535, 0.0003063596, 0,
  0, 0, 0.0003063596, 0.00161393, 0.002611525, 0.002611525, 0.00161393, 
    0.0003063596, 0, 0,
  0, 0, 0, 0.0004326566, 0.0007000027, 0.0007000027, 0.0004326566, 0, 0, 0,
  0, 0, 0, 0.0003493234, 0.0005684707, 0.0005684707, 0.0003493234, 0, 0, 0,
  0, 0, 0.0002173396, 0.001303148, 0.002120834, 0.002120834, 0.001303148, 
    0.0002173396, 0, 0,
  0, 0.0002173396, 0.007451856, 0.006906761, 0.00616609, 0.00616609, 
    0.006906761, 0.007451856, 0.0002173396, 0,
  0.0003493234, 0.001303148, 0.006906761, 0.003873749, 0.001350252, 
    0.001350252, 0.003873749, 0.006906761, 0.001303148, 0.0003493234,
  0.0005684707, 0.002120834, 0.00616609, 0.001350252, 8.674125e-05, 
    8.674125e-05, 0.001350252, 0.00616609, 0.002120834, 0.0005684707,
  0.0005684707, 0.002120834, 0.00616609, 0.001350252, 8.674125e-05, 
    8.674125e-05, 0.001350252, 0.00616609, 0.002120834, 0.0005684707,
  0.0003493234, 0.001303148, 0.006906761, 0.003873749, 0.001350252, 
    0.001350252, 0.003873749, 0.006906761, 0.001303148, 0.0003493234,
  0, 0.0002173396, 0.007451856, 0.006906761, 0.00616609, 0.00616609, 
    0.006906761, 0.007451856, 0.0002173396, 0,
  0, 0, 0.0002173396, 0.001303148, 0.002120834, 0.002120834, 0.001303148, 
    0.0002173396, 0, 0,
  0, 0, 0, 0.0003493234, 0.0005684707, 0.0005684707, 0.0003493234, 0, 0, 0,
  0, 0, 0, 0.0002606724, 0.0004258991, 0.0004258991, 0.0002606724, 0, 0, 0,
  0, 0, 0.0001459482, 0.0009725092, 0.001589012, 0.001589012, 0.0009725092, 
    0.0001459482, 0, 0,
  0, 0.0001459482, 0.005637544, 0.005234025, 0.00467806, 0.00467806, 
    0.005234025, 0.005637544, 0.0001459482, 0,
  0.0002606724, 0.0009725092, 0.005234025, 0.002913182, 0.001005295, 
    0.001005295, 0.002913182, 0.005234025, 0.0009725092, 0.0002606724,
  0.0004258991, 0.001589012, 0.00467806, 0.001005295, 6.351428e-05, 
    6.351428e-05, 0.001005295, 0.00467806, 0.001589012, 0.0004258991,
  0.0004258991, 0.001589012, 0.00467806, 0.001005295, 6.351428e-05, 
    6.351428e-05, 0.001005295, 0.00467806, 0.001589012, 0.0004258991,
  0.0002606724, 0.0009725092, 0.005234025, 0.002913182, 0.001005295, 
    0.001005295, 0.002913182, 0.005234025, 0.0009725092, 0.0002606724,
  0, 0.0001459482, 0.005637544, 0.005234025, 0.00467806, 0.00467806, 
    0.005234025, 0.005637544, 0.0001459482, 0,
  0, 0, 0.0001459482, 0.0009725092, 0.001589012, 0.001589012, 0.0009725092, 
    0.0001459482, 0, 0,
  0, 0, 0, 0.0002606724, 0.0004258991, 0.0004258991, 0.0002606724, 0, 0, 0,
  0, 0, 0, 0.0001712833, 0.0002805443, 0.0002805443, 0.0001712833, 0, 0, 0,
  0, 0, 8.849078e-05, 0.0006390744, 0.001046777, 0.001046777, 0.0006390744, 
    8.849078e-05, 0, 0,
  0, 8.849078e-05, 0.003750738, 0.00348681, 0.003119645, 0.003119645, 
    0.00348681, 0.003750738, 8.849078e-05, 0,
  0.0001712833, 0.0006390744, 0.00348681, 0.001927426, 0.0006600972, 
    0.0006600972, 0.001927426, 0.00348681, 0.0006390744, 0.0001712833,
  0.0002805443, 0.001046777, 0.003119645, 0.0006600972, 4.144524e-05, 
    4.144524e-05, 0.0006600972, 0.003119645, 0.001046777, 0.0002805443,
  0.0002805443, 0.001046777, 0.003119645, 0.0006600972, 4.144524e-05, 
    4.144524e-05, 0.0006600972, 0.003119645, 0.001046777, 0.0002805443,
  0.0001712833, 0.0006390744, 0.00348681, 0.001927426, 0.0006600972, 
    0.0006600972, 0.001927426, 0.00348681, 0.0006390744, 0.0001712833,
  0, 8.849078e-05, 0.003750738, 0.00348681, 0.003119645, 0.003119645, 
    0.00348681, 0.003750738, 8.849078e-05, 0,
  0, 0, 8.849078e-05, 0.0006390744, 0.001046777, 0.001046777, 0.0006390744, 
    8.849078e-05, 0, 0,
  0, 0, 0, 0.0001712833, 0.0002805443, 0.0002805443, 0.0001712833, 0, 0, 0,
  0, 0, 0, 8.390821e-05, 0.0001376783, 0.0001376783, 8.390821e-05, 0, 0, 0,
  0, 0, 4.070004e-05, 0.0003131028, 0.0005137604, 0.0005137604, 0.0003131028, 
    4.070004e-05, 0, 0,
  0, 4.070004e-05, 0.00186055, 0.001732983, 0.001552684, 0.001552684, 
    0.001732983, 0.00186055, 4.070004e-05, 0,
  8.390821e-05, 0.0003131028, 0.001732983, 0.0009527217, 0.0003241294, 
    0.0003241294, 0.0009527217, 0.001732983, 0.0003131028, 8.390821e-05,
  0.0001376783, 0.0005137604, 0.001552684, 0.0003241294, 2.035775e-05, 
    2.035775e-05, 0.0003241294, 0.001552684, 0.0005137604, 0.0001376783,
  0.0001376783, 0.0005137604, 0.001552684, 0.0003241294, 2.035775e-05, 
    2.035775e-05, 0.0003241294, 0.001552684, 0.0005137604, 0.0001376783,
  8.390821e-05, 0.0003131028, 0.001732983, 0.0009527217, 0.0003241294, 
    0.0003241294, 0.0009527217, 0.001732983, 0.0003131028, 8.390821e-05,
  0, 4.070004e-05, 0.00186055, 0.001732983, 0.001552684, 0.001552684, 
    0.001732983, 0.00186055, 4.070004e-05, 0,
  0, 0, 4.070004e-05, 0.0003131028, 0.0005137604, 0.0005137604, 0.0003131028, 
    4.070004e-05, 0, 0,
  0, 0, 0, 8.390821e-05, 0.0001376783, 0.0001376783, 8.390821e-05, 0, 0, 0,
  0, 0, 0, 5.844771e-09, 7.009599e-09, 7.009599e-09, 5.844771e-09, 0, 0, 0,
  0, 0, 1.757822e-08, 2.418835e-08, 2.870435e-08, 2.870435e-08, 2.418835e-08, 
    1.757822e-08, 0, 0,
  0, 1.757822e-08, 3.317751e-08, 2.910274e-08, 2.583801e-08, 2.583801e-08, 
    2.910274e-08, 3.317751e-08, 1.757822e-08, 0,
  5.844771e-09, 2.418835e-08, 2.910274e-08, 2.178858e-08, 1.614761e-08, 
    1.614761e-08, 2.178858e-08, 2.910274e-08, 2.418835e-08, 5.844771e-09,
  7.009599e-09, 2.870435e-08, 2.583801e-08, 1.614761e-08, 8.26189e-09, 
    8.26189e-09, 1.614761e-08, 2.583801e-08, 2.870435e-08, 7.009599e-09,
  7.009599e-09, 2.870435e-08, 2.583801e-08, 1.614761e-08, 8.26189e-09, 
    8.26189e-09, 1.614761e-08, 2.583801e-08, 2.870435e-08, 7.009599e-09,
  5.844771e-09, 2.418835e-08, 2.910274e-08, 2.178858e-08, 1.614761e-08, 
    1.614761e-08, 2.178858e-08, 2.910274e-08, 2.418835e-08, 5.844771e-09,
  0, 1.757822e-08, 3.317751e-08, 2.910274e-08, 2.583801e-08, 2.583801e-08, 
    2.910274e-08, 3.317751e-08, 1.757822e-08, 0,
  0, 0, 1.757822e-08, 2.418835e-08, 2.870435e-08, 2.870435e-08, 2.418835e-08, 
    1.757822e-08, 0, 0,
  0, 0, 0, 5.844771e-09, 7.009599e-09, 7.009599e-09, 5.844771e-09, 0, 0, 0,
  0, 0, 0, 0.0006069986, 0.00093498, 0.00093498, 0.0006069986, 0, 0, 0,
  0, 0, 0.0007784671, 0.002264374, 0.003496286, 0.003496286, 0.002264374, 
    0.0007784671, 0, 0,
  0, 0.0007784671, 0.01173998, 0.01082779, 0.009718124, 0.009718124, 
    0.01082779, 0.01173998, 0.0007784671, 0,
  0.0006069986, 0.002264374, 0.01082779, 0.006453543, 0.002536954, 
    0.002536954, 0.006453543, 0.01082779, 0.002264374, 0.0006069986,
  0.00093498, 0.003496286, 0.009718124, 0.002536954, 0.0002054527, 
    0.0002054527, 0.002536954, 0.009718124, 0.003496286, 0.00093498,
  0.00093498, 0.003496286, 0.009718124, 0.002536954, 0.0002054527, 
    0.0002054527, 0.002536954, 0.009718124, 0.003496286, 0.00093498,
  0.0006069986, 0.002264374, 0.01082779, 0.006453543, 0.002536954, 
    0.002536954, 0.006453543, 0.01082779, 0.002264374, 0.0006069986,
  0, 0.0007784671, 0.01173998, 0.01082779, 0.009718124, 0.009718124, 
    0.01082779, 0.01173998, 0.0007784671, 0,
  0, 0, 0.0007784671, 0.002264374, 0.003496286, 0.003496286, 0.002264374, 
    0.0007784671, 0, 0,
  0, 0, 0, 0.0006069986, 0.00093498, 0.00093498, 0.0006069986, 0, 0, 0,
  0, 0, 0, 0.0005942544, 0.0009234856, 0.0009234856, 0.0005942544, 0, 0, 0,
  0, 0, 0.0007008232, 0.002216507, 0.003448871, 0.003448871, 0.002216507, 
    0.0007008232, 0, 0,
  0, 0.0007008232, 0.0116403, 0.01070889, 0.009588439, 0.009588439, 
    0.01070889, 0.0116403, 0.0007008232, 0,
  0.0005942544, 0.002216507, 0.01070889, 0.006344839, 0.002455897, 
    0.002455897, 0.006344839, 0.01070889, 0.002216507, 0.0005942544,
  0.0009234856, 0.003448871, 0.009588439, 0.002455897, 0.0001934233, 
    0.0001934233, 0.002455897, 0.009588439, 0.003448871, 0.0009234856,
  0.0009234856, 0.003448871, 0.009588439, 0.002455897, 0.0001934233, 
    0.0001934233, 0.002455897, 0.009588439, 0.003448871, 0.0009234856,
  0.0005942544, 0.002216507, 0.01070889, 0.006344839, 0.002455897, 
    0.002455897, 0.006344839, 0.01070889, 0.002216507, 0.0005942544,
  0, 0.0007008232, 0.0116403, 0.01070889, 0.009588439, 0.009588439, 
    0.01070889, 0.0116403, 0.0007008232, 0,
  0, 0, 0.0007008232, 0.002216507, 0.003448871, 0.003448871, 0.002216507, 
    0.0007008232, 0, 0,
  0, 0, 0, 0.0005942544, 0.0009234856, 0.0009234856, 0.0005942544, 0, 0, 0,
  0, 0, 0, 0.0005617622, 0.0008875804, 0.0008875804, 0.0005617622, 0, 0, 0,
  0, 0, 0.0005628115, 0.002095515, 0.003312497, 0.003312497, 0.002095515, 
    0.0005628115, 0, 0,
  0, 0.0005628115, 0.01126161, 0.01033729, 0.009212223, 0.009212223, 
    0.01033729, 0.01126161, 0.0005628115, 0,
  0.0005617622, 0.002095515, 0.01033729, 0.006014444, 0.002253723, 
    0.002253723, 0.006014444, 0.01033729, 0.002095515, 0.0005617622,
  0.0008875804, 0.003312497, 0.009212223, 0.002253723, 0.000169539, 
    0.000169539, 0.002253723, 0.009212223, 0.003312497, 0.0008875804,
  0.0008875804, 0.003312497, 0.009212223, 0.002253723, 0.000169539, 
    0.000169539, 0.002253723, 0.009212223, 0.003312497, 0.0008875804,
  0.0005617622, 0.002095515, 0.01033729, 0.006014444, 0.002253723, 
    0.002253723, 0.006014444, 0.01033729, 0.002095515, 0.0005617622,
  0, 0.0005628115, 0.01126161, 0.01033729, 0.009212223, 0.009212223, 
    0.01033729, 0.01126161, 0.0005628115, 0,
  0, 0, 0.0005628115, 0.002095515, 0.003312497, 0.003312497, 0.002095515, 
    0.0005628115, 0, 0,
  0, 0, 0, 0.0005617622, 0.0008875804, 0.0008875804, 0.0005617622, 0, 0, 0,
  0, 0, 0, 0.0005082712, 0.0008128783, 0.0008128783, 0.0005082712, 0, 0, 0,
  0, 0, 0.0004322867, 0.001895953, 0.003032888, 0.003032888, 0.001895953, 
    0.0004322867, 0, 0,
  0, 0.0004322867, 0.01040767, 0.009564335, 0.008505442, 0.008505442, 
    0.009564335, 0.01040767, 0.0004322867, 0,
  0.0005082712, 0.001895953, 0.009564335, 0.005476218, 0.00199077, 
    0.00199077, 0.005476218, 0.009564335, 0.001895953, 0.0005082712,
  0.0008128783, 0.003032888, 0.008505442, 0.00199077, 0.0001412429, 
    0.0001412429, 0.00199077, 0.008505442, 0.003032888, 0.0008128783,
  0.0008128783, 0.003032888, 0.008505442, 0.00199077, 0.0001412429, 
    0.0001412429, 0.00199077, 0.008505442, 0.003032888, 0.0008128783,
  0.0005082712, 0.001895953, 0.009564335, 0.005476218, 0.00199077, 
    0.00199077, 0.005476218, 0.009564335, 0.001895953, 0.0005082712,
  0, 0.0004322867, 0.01040767, 0.009564335, 0.008505442, 0.008505442, 
    0.009564335, 0.01040767, 0.0004322867, 0,
  0, 0, 0.0004322867, 0.001895953, 0.003032888, 0.003032888, 0.001895953, 
    0.0004322867, 0, 0,
  0, 0, 0, 0.0005082712, 0.0008128783, 0.0008128783, 0.0005082712, 0, 0, 0,
  0, 0, 0, 0.0004361948, 0.0007032796, 0.0007032796, 0.0004361948, 0, 0, 0,
  0, 0, 0.0003210134, 0.00162713, 0.002623765, 0.002623765, 0.00162713, 
    0.0003210134, 0, 0,
  0, 0.0003210134, 0.009096134, 0.008377466, 0.007451397, 0.007451397, 
    0.008377466, 0.009096134, 0.0003210134, 0,
  0.0004361948, 0.00162713, 0.008377466, 0.004740235, 0.001687256, 
    0.001687256, 0.004740235, 0.008377466, 0.00162713, 0.0004361948,
  0.0007032796, 0.002623765, 0.007451397, 0.001687256, 0.0001137157, 
    0.0001137157, 0.001687256, 0.007451397, 0.002623765, 0.0007032796,
  0.0007032796, 0.002623765, 0.007451397, 0.001687256, 0.0001137157, 
    0.0001137157, 0.001687256, 0.007451397, 0.002623765, 0.0007032796,
  0.0004361948, 0.00162713, 0.008377466, 0.004740235, 0.001687256, 
    0.001687256, 0.004740235, 0.008377466, 0.00162713, 0.0004361948,
  0, 0.0003210134, 0.009096134, 0.008377466, 0.007451397, 0.007451397, 
    0.008377466, 0.009096134, 0.0003210134, 0,
  0, 0, 0.0003210134, 0.00162713, 0.002623765, 0.002623765, 0.00162713, 
    0.0003210134, 0, 0,
  0, 0, 0, 0.0004361948, 0.0007032796, 0.0007032796, 0.0004361948, 0, 0, 0,
  0, 0, 0, 0.0003522951, 0.0005712211, 0.0005712211, 0.0003522951, 0, 0, 0,
  0, 0, 0.0002289628, 0.001314233, 0.002131102, 0.002131102, 0.001314233, 
    0.0002289628, 0, 0,
  0, 0.0002289628, 0.007463273, 0.006887882, 0.006132556, 0.006132556, 
    0.006887882, 0.007463273, 0.0002289628, 0,
  0.0003522951, 0.001314233, 0.006887882, 0.003861439, 0.001355211, 
    0.001355211, 0.003861439, 0.006887882, 0.001314233, 0.0003522951,
  0.0005712211, 0.002131102, 0.006132556, 0.001355211, 8.841011e-05, 
    8.841011e-05, 0.001355211, 0.006132556, 0.002131102, 0.0005712211,
  0.0005712211, 0.002131102, 0.006132556, 0.001355211, 8.841011e-05, 
    8.841011e-05, 0.001355211, 0.006132556, 0.002131102, 0.0005712211,
  0.0003522951, 0.001314233, 0.006887882, 0.003861439, 0.001355211, 
    0.001355211, 0.003861439, 0.006887882, 0.001314233, 0.0003522951,
  0, 0.0002289628, 0.007463273, 0.006887882, 0.006132556, 0.006132556, 
    0.006887882, 0.007463273, 0.0002289628, 0,
  0, 0, 0.0002289628, 0.001314233, 0.002131102, 0.002131102, 0.001314233, 
    0.0002289628, 0, 0,
  0, 0, 0, 0.0003522951, 0.0005712211, 0.0005712211, 0.0003522951, 0, 0, 0,
  0, 0, 0, 0.0002629973, 0.0004280503, 0.0004280503, 0.0002629973, 0, 0, 0,
  0, 0, 0.0001544167, 0.0009811802, 0.001597041, 0.001597041, 0.0009811802, 
    0.0001544167, 0, 0,
  0, 0.0001544167, 0.005649096, 0.005221925, 0.004654344, 0.004654344, 
    0.005221925, 0.005649096, 0.0001544167, 0,
  0.0002629973, 0.0009811802, 0.005221925, 0.002904604, 0.001009367, 
    0.001009367, 0.002904604, 0.005221925, 0.0009811802, 0.0002629973,
  0.0004280503, 0.001597041, 0.004654344, 0.001009367, 6.476569e-05, 
    6.476569e-05, 0.001009367, 0.004654344, 0.001597041, 0.0004280503,
  0.0004280503, 0.001597041, 0.004654344, 0.001009367, 6.476569e-05, 
    6.476569e-05, 0.001009367, 0.004654344, 0.001597041, 0.0004280503,
  0.0002629973, 0.0009811802, 0.005221925, 0.002904604, 0.001009367, 
    0.001009367, 0.002904604, 0.005221925, 0.0009811802, 0.0002629973,
  0, 0.0001544167, 0.005649096, 0.005221925, 0.004654344, 0.004654344, 
    0.005221925, 0.005649096, 0.0001544167, 0,
  0, 0, 0.0001544167, 0.0009811802, 0.001597041, 0.001597041, 0.0009811802, 
    0.0001544167, 0, 0,
  0, 0, 0, 0.0002629973, 0.0004280503, 0.0004280503, 0.0002629973, 0, 0, 0,
  0, 0, 0, 0.0001728918, 0.0002820509, 0.0002820509, 0.0001728918, 0, 0, 0,
  0, 0, 9.381691e-05, 0.0006450738, 0.001052398, 0.001052398, 0.0006450738, 
    9.381691e-05, 0, 0,
  0, 9.381691e-05, 0.003761029, 0.003481176, 0.003105961, 0.003105961, 
    0.003481176, 0.003761029, 9.381691e-05, 0,
  0.0001728918, 0.0006450738, 0.003481176, 0.001922795, 0.0006631501, 
    0.0006631501, 0.001922795, 0.003481176, 0.0006450738, 0.0001728918,
  0.0002820509, 0.001052398, 0.003105961, 0.0006631501, 4.229241e-05, 
    4.229241e-05, 0.0006631501, 0.003105961, 0.001052398, 0.0002820509,
  0.0002820509, 0.001052398, 0.003105961, 0.0006631501, 4.229241e-05, 
    4.229241e-05, 0.0006631501, 0.003105961, 0.001052398, 0.0002820509,
  0.0001728918, 0.0006450738, 0.003481176, 0.001922795, 0.0006631501, 
    0.0006631501, 0.001922795, 0.003481176, 0.0006450738, 0.0001728918,
  0, 9.381691e-05, 0.003761029, 0.003481176, 0.003105961, 0.003105961, 
    0.003481176, 0.003761029, 9.381691e-05, 0,
  0, 0, 9.381691e-05, 0.0006450738, 0.001052398, 0.001052398, 0.0006450738, 
    9.381691e-05, 0, 0,
  0, 0, 0, 0.0001728918, 0.0002820509, 0.0002820509, 0.0001728918, 0, 0, 0,
  0, 0, 0, 8.472346e-05, 0.0001384727, 0.0001384727, 8.472346e-05, 0, 0, 0,
  0, 0, 4.305005e-05, 0.0003161442, 0.0005167247, 0.0005167247, 0.0003161442, 
    4.305005e-05, 0, 0,
  0, 4.305005e-05, 0.001866988, 0.001731893, 0.001547656, 0.001547656, 
    0.001731893, 0.001866988, 4.305005e-05, 0,
  8.472346e-05, 0.0003161442, 0.001731893, 0.0009515861, 0.0003259962, 
    0.0003259962, 0.0009515861, 0.001731893, 0.0003161442, 8.472346e-05,
  0.0001384727, 0.0005167247, 0.001547656, 0.0003259962, 2.079849e-05, 
    2.079849e-05, 0.0003259962, 0.001547656, 0.0005167247, 0.0001384727,
  0.0001384727, 0.0005167247, 0.001547656, 0.0003259962, 2.079849e-05, 
    2.079849e-05, 0.0003259962, 0.001547656, 0.0005167247, 0.0001384727,
  8.472346e-05, 0.0003161442, 0.001731893, 0.0009515861, 0.0003259962, 
    0.0003259962, 0.0009515861, 0.001731893, 0.0003161442, 8.472346e-05,
  0, 4.305005e-05, 0.001866988, 0.001731893, 0.001547656, 0.001547656, 
    0.001731893, 0.001866988, 4.305005e-05, 0,
  0, 0, 4.305005e-05, 0.0003161442, 0.0005167247, 0.0005167247, 0.0003161442, 
    4.305005e-05, 0, 0,
  0, 0, 0, 8.472346e-05, 0.0001384727, 0.0001384727, 8.472346e-05, 0, 0, 0,
  0, 0, 0, 5.848141e-09, 7.010175e-09, 7.010175e-09, 5.848141e-09, 0, 0, 0,
  0, 0, 1.76082e-08, 2.421836e-08, 2.872793e-08, 2.872793e-08, 2.421836e-08, 
    1.76082e-08, 0, 0,
  0, 1.76082e-08, 3.316813e-08, 2.905329e-08, 2.576806e-08, 2.576806e-08, 
    2.905329e-08, 3.316813e-08, 1.76082e-08, 0,
  5.848141e-09, 2.421836e-08, 2.905329e-08, 2.176385e-08, 1.61552e-08, 
    1.61552e-08, 2.176385e-08, 2.905329e-08, 2.421836e-08, 5.848141e-09,
  7.010175e-09, 2.872793e-08, 2.576806e-08, 1.61552e-08, 8.291257e-09, 
    8.291257e-09, 1.61552e-08, 2.576806e-08, 2.872793e-08, 7.010175e-09,
  7.010175e-09, 2.872793e-08, 2.576806e-08, 1.61552e-08, 8.291257e-09, 
    8.291257e-09, 1.61552e-08, 2.576806e-08, 2.872793e-08, 7.010175e-09,
  5.848141e-09, 2.421836e-08, 2.905329e-08, 2.176385e-08, 1.61552e-08, 
    1.61552e-08, 2.176385e-08, 2.905329e-08, 2.421836e-08, 5.848141e-09,
  0, 1.76082e-08, 3.316813e-08, 2.905329e-08, 2.576806e-08, 2.576806e-08, 
    2.905329e-08, 3.316813e-08, 1.76082e-08, 0,
  0, 0, 1.76082e-08, 2.421836e-08, 2.872793e-08, 2.872793e-08, 2.421836e-08, 
    1.76082e-08, 0, 0,
  0, 0, 0, 5.848141e-09, 7.010175e-09, 7.010175e-09, 5.848141e-09, 0, 0, 0,
  0, 0, 0, 0.0006112515, 0.0009389082, 0.0009389082, 0.0006112515, 0, 0, 0,
  0, 0, 0.0007980737, 0.002280353, 0.003511114, 0.003511114, 0.002280353, 
    0.0007980737, 0, 0,
  0, 0.0007980737, 0.01174879, 0.0107924, 0.009659738, 0.009659738, 
    0.0107924, 0.01174879, 0.0007980737, 0,
  0.0006112515, 0.002280353, 0.0107924, 0.00643165, 0.002542179, 0.002542179, 
    0.00643165, 0.0107924, 0.002280353, 0.0006112515,
  0.0009389082, 0.003511114, 0.009659738, 0.002542179, 0.0002090917, 
    0.0002090917, 0.002542179, 0.009659738, 0.003511114, 0.0009389082,
  0.0009389082, 0.003511114, 0.009659738, 0.002542179, 0.0002090917, 
    0.0002090917, 0.002542179, 0.009659738, 0.003511114, 0.0009389082,
  0.0006112515, 0.002280353, 0.0107924, 0.00643165, 0.002542179, 0.002542179, 
    0.00643165, 0.0107924, 0.002280353, 0.0006112515,
  0, 0.0007980737, 0.01174879, 0.0107924, 0.009659738, 0.009659738, 
    0.0107924, 0.01174879, 0.0007980737, 0,
  0, 0, 0.0007980737, 0.002280353, 0.003511114, 0.003511114, 0.002280353, 
    0.0007980737, 0, 0,
  0, 0, 0, 0.0006112515, 0.0009389082, 0.0009389082, 0.0006112515, 0, 0, 0,
  0, 0, 0, 0.0005985127, 0.0009274351, 0.0009274351, 0.0005985127, 0, 0, 0,
  0, 0, 0.0007204616, 0.002232448, 0.0034637, 0.0034637, 0.002232448, 
    0.0007204616, 0, 0,
  0, 0.0007204616, 0.01164908, 0.01067409, 0.009531437, 0.009531437, 
    0.01067409, 0.01164908, 0.0007204616, 0,
  0.0005985127, 0.002232448, 0.01067409, 0.00632325, 0.002461222, 
    0.002461222, 0.00632325, 0.01067409, 0.002232448, 0.0005985127,
  0.0009274351, 0.0034637, 0.009531437, 0.002461222, 0.0001968937, 
    0.0001968937, 0.002461222, 0.009531437, 0.0034637, 0.0009274351,
  0.0009274351, 0.0034637, 0.009531437, 0.002461222, 0.0001968937, 
    0.0001968937, 0.002461222, 0.009531437, 0.0034637, 0.0009274351,
  0.0005985127, 0.002232448, 0.01067409, 0.00632325, 0.002461222, 
    0.002461222, 0.00632325, 0.01067409, 0.002232448, 0.0005985127,
  0, 0.0007204616, 0.01164908, 0.01067409, 0.009531437, 0.009531437, 
    0.01067409, 0.01164908, 0.0007204616, 0,
  0, 0, 0.0007204616, 0.002232448, 0.0034637, 0.0034637, 0.002232448, 
    0.0007204616, 0, 0,
  0, 0, 0, 0.0005985127, 0.0009274351, 0.0009274351, 0.0005985127, 0, 0, 0,
  0, 0, 0, 0.0005659737, 0.0008914738, 0.0008914738, 0.0005659737, 0, 0, 0,
  0, 0, 0.0005818107, 0.002111247, 0.003327071, 0.003327071, 0.002111247, 
    0.0005818107, 0, 0,
  0, 0.0005818107, 0.0112707, 0.0103041, 0.009158306, 0.009158306, 0.0103041, 
    0.0112707, 0.0005818107, 0,
  0.0005659737, 0.002111247, 0.0103041, 0.005994077, 0.002259386, 
    0.002259386, 0.005994077, 0.0103041, 0.002111247, 0.0005659737,
  0.0008914738, 0.003327071, 0.009158306, 0.002259386, 0.0001725932, 
    0.0001725932, 0.002259386, 0.009158306, 0.003327071, 0.0008914738,
  0.0008914738, 0.003327071, 0.009158306, 0.002259386, 0.0001725932, 
    0.0001725932, 0.002259386, 0.009158306, 0.003327071, 0.0008914738,
  0.0005659737, 0.002111247, 0.0103041, 0.005994077, 0.002259386, 
    0.002259386, 0.005994077, 0.0103041, 0.002111247, 0.0005659737,
  0, 0.0005818107, 0.0112707, 0.0103041, 0.009158306, 0.009158306, 0.0103041, 
    0.0112707, 0.0005818107, 0,
  0, 0, 0.0005818107, 0.002111247, 0.003327071, 0.003327071, 0.002111247, 
    0.0005818107, 0, 0,
  0, 0, 0, 0.0005659737, 0.0008914738, 0.0008914738, 0.0005659737, 0, 0, 0,
  0, 0, 0, 0.0005122339, 0.0008165314, 0.0008165314, 0.0005122339, 0, 0, 0,
  0, 0, 0.0004496239, 0.001910743, 0.003046544, 0.003046544, 0.001910743, 
    0.0004496239, 0, 0,
  0, 0.0004496239, 0.0104174, 0.009534373, 0.008456479, 0.008456479, 
    0.009534373, 0.0104174, 0.0004496239, 0,
  0.0005122339, 0.001910743, 0.009534373, 0.0054579, 0.001996574, 
    0.001996574, 0.0054579, 0.009534373, 0.001910743, 0.0005122339,
  0.0008165314, 0.003046544, 0.008456479, 0.001996574, 0.0001438155, 
    0.0001438155, 0.001996574, 0.008456479, 0.003046544, 0.0008165314,
  0.0008165314, 0.003046544, 0.008456479, 0.001996574, 0.0001438155, 
    0.0001438155, 0.001996574, 0.008456479, 0.003046544, 0.0008165314,
  0.0005122339, 0.001910743, 0.009534373, 0.0054579, 0.001996574, 
    0.001996574, 0.0054579, 0.009534373, 0.001910743, 0.0005122339,
  0, 0.0004496239, 0.0104174, 0.009534373, 0.008456479, 0.008456479, 
    0.009534373, 0.0104174, 0.0004496239, 0,
  0, 0, 0.0004496239, 0.001910743, 0.003046544, 0.003046544, 0.001910743, 
    0.0004496239, 0, 0,
  0, 0, 0, 0.0005122339, 0.0008165314, 0.0008165314, 0.0005122339, 0, 0, 0,
  0, 0, 0, 0.0004397197, 0.000706529, 0.000706529, 0.0004397197, 0, 0, 0,
  0, 0, 0.0003358313, 0.00164028, 0.002635903, 0.002635903, 0.00164028, 
    0.0003358313, 0, 0,
  0, 0.0003358313, 0.009106624, 0.008352441, 0.007409481, 0.007409481, 
    0.008352441, 0.009106624, 0.0003358313, 0,
  0.0004397197, 0.00164028, 0.008352441, 0.0047247, 0.001692774, 0.001692774, 
    0.0047247, 0.008352441, 0.00164028, 0.0004397197,
  0.000706529, 0.002635903, 0.007409481, 0.001692774, 0.0001158285, 
    0.0001158285, 0.001692774, 0.007409481, 0.002635903, 0.000706529,
  0.000706529, 0.002635903, 0.007409481, 0.001692774, 0.0001158285, 
    0.0001158285, 0.001692774, 0.007409481, 0.002635903, 0.000706529,
  0.0004397197, 0.00164028, 0.008352441, 0.0047247, 0.001692774, 0.001692774, 
    0.0047247, 0.008352441, 0.00164028, 0.0004397197,
  0, 0.0003358313, 0.009106624, 0.008352441, 0.007409481, 0.007409481, 
    0.008352441, 0.009106624, 0.0003358313, 0,
  0, 0, 0.0003358313, 0.00164028, 0.002635903, 0.002635903, 0.00164028, 
    0.0003358313, 0, 0,
  0, 0, 0, 0.0004397197, 0.000706529, 0.000706529, 0.0004397197, 0, 0, 0,
  0, 0, 0, 0.0003552552, 0.0005739492, 0.0005739492, 0.0003552552, 0, 0, 0,
  0, 0, 0.0002408023, 0.001325274, 0.002141288, 0.002141288, 0.001325274, 
    0.0002408023, 0, 0,
  0, 0.0002408023, 0.007474388, 0.006869011, 0.006099347, 0.006099347, 
    0.006869011, 0.007474388, 0.0002408023, 0,
  0.0003552552, 0.001325274, 0.006869011, 0.003849247, 0.001360088, 
    0.001360088, 0.003849247, 0.006869011, 0.001325274, 0.0003552552,
  0.0005739492, 0.002141288, 0.006099347, 0.001360088, 9.00874e-05, 
    9.00874e-05, 0.001360088, 0.006099347, 0.002141288, 0.0005739492,
  0.0005739492, 0.002141288, 0.006099347, 0.001360088, 9.00874e-05, 
    9.00874e-05, 0.001360088, 0.006099347, 0.002141288, 0.0005739492,
  0.0003552552, 0.001325274, 0.006869011, 0.003849247, 0.001360088, 
    0.001360088, 0.003849247, 0.006869011, 0.001325274, 0.0003552552,
  0, 0.0002408023, 0.007474388, 0.006869011, 0.006099347, 0.006099347, 
    0.006869011, 0.007474388, 0.0002408023, 0,
  0, 0, 0.0002408023, 0.001325274, 0.002141288, 0.002141288, 0.001325274, 
    0.0002408023, 0, 0,
  0, 0, 0, 0.0003552552, 0.0005739492, 0.0005739492, 0.0003552552, 0, 0, 0,
  0, 0, 0, 0.0002653098, 0.0004301848, 0.0004301848, 0.0002653098, 0, 0, 0,
  0, 0, 0.0001631102, 0.0009898049, 0.001605008, 0.001605008, 0.0009898049, 
    0.0001631102, 0, 0,
  0, 0.0001631102, 0.005660271, 0.005209757, 0.004630838, 0.004630838, 
    0.005209757, 0.005660271, 0.0001631102, 0,
  0.0002653098, 0.0009898049, 0.005209757, 0.002896127, 0.001013378, 
    0.001013378, 0.002896127, 0.005209757, 0.0009898049, 0.0002653098,
  0.0004301848, 0.001605008, 0.004630838, 0.001013378, 6.602427e-05, 
    6.602427e-05, 0.001013378, 0.004630838, 0.001605008, 0.0004301848,
  0.0004301848, 0.001605008, 0.004630838, 0.001013378, 6.602427e-05, 
    6.602427e-05, 0.001013378, 0.004630838, 0.001605008, 0.0004301848,
  0.0002653098, 0.0009898049, 0.005209757, 0.002896127, 0.001013378, 
    0.001013378, 0.002896127, 0.005209757, 0.0009898049, 0.0002653098,
  0, 0.0001631102, 0.005660271, 0.005209757, 0.004630838, 0.004630838, 
    0.005209757, 0.005660271, 0.0001631102, 0,
  0, 0, 0.0001631102, 0.0009898049, 0.001605008, 0.001605008, 0.0009898049, 
    0.0001631102, 0, 0,
  0, 0, 0, 0.0002653098, 0.0004301848, 0.0004301848, 0.0002653098, 0, 0, 0,
  0, 0, 0, 0.0001744839, 0.0002835433, 0.0002835433, 0.0001744839, 0, 0, 0,
  0, 0, 9.931539e-05, 0.0006510119, 0.001057967, 0.001057967, 0.0006510119, 
    9.931539e-05, 0, 0,
  0, 9.931539e-05, 0.003770805, 0.003475333, 0.003092316, 0.003092316, 
    0.003475333, 0.003770805, 9.931539e-05, 0,
  0.0001744839, 0.0006510119, 0.003475333, 0.001918233, 0.0006661618, 
    0.0006661618, 0.001918233, 0.003475333, 0.0006510119, 0.0001744839,
  0.0002835433, 0.001057967, 0.003092316, 0.0006661618, 4.314424e-05, 
    4.314424e-05, 0.0006661618, 0.003092316, 0.001057967, 0.0002835433,
  0.0002835433, 0.001057967, 0.003092316, 0.0006661618, 4.314424e-05, 
    4.314424e-05, 0.0006661618, 0.003092316, 0.001057967, 0.0002835433,
  0.0001744839, 0.0006510119, 0.003475333, 0.001918233, 0.0006661618, 
    0.0006661618, 0.001918233, 0.003475333, 0.0006510119, 0.0001744839,
  0, 9.931539e-05, 0.003770805, 0.003475333, 0.003092316, 0.003092316, 
    0.003475333, 0.003770805, 9.931539e-05, 0,
  0, 0, 9.931539e-05, 0.0006510119, 0.001057967, 0.001057967, 0.0006510119, 
    9.931539e-05, 0, 0,
  0, 0, 0, 0.0001744839, 0.0002835433, 0.0002835433, 0.0001744839, 0, 0, 0,
  0, 0, 0, 8.552483e-05, 0.0001392532, 0.0001392532, 8.552483e-05, 0, 0, 0,
  0, 0, 4.550071e-05, 0.0003191338, 0.000519637, 0.000519637, 0.0003191338, 
    4.550071e-05, 0, 0,
  0, 4.550071e-05, 0.001872948, 0.001730472, 0.001542442, 0.001542442, 
    0.001730472, 0.001872948, 4.550071e-05, 0,
  8.552483e-05, 0.0003191338, 0.001730472, 0.0009503962, 0.0003278269, 
    0.0003278269, 0.0009503962, 0.001730472, 0.0003191338, 8.552483e-05,
  0.0001392532, 0.000519637, 0.001542442, 0.0003278269, 2.123982e-05, 
    2.123982e-05, 0.0003278269, 0.001542442, 0.000519637, 0.0001392532,
  0.0001392532, 0.000519637, 0.001542442, 0.0003278269, 2.123982e-05, 
    2.123982e-05, 0.0003278269, 0.001542442, 0.000519637, 0.0001392532,
  8.552483e-05, 0.0003191338, 0.001730472, 0.0009503962, 0.0003278269, 
    0.0003278269, 0.0009503962, 0.001730472, 0.0003191338, 8.552483e-05,
  0, 4.550071e-05, 0.001872948, 0.001730472, 0.001542442, 0.001542442, 
    0.001730472, 0.001872948, 4.550071e-05, 0,
  0, 0, 4.550071e-05, 0.0003191338, 0.000519637, 0.000519637, 0.0003191338, 
    4.550071e-05, 0, 0,
  0, 0, 0, 8.552483e-05, 0.0001392532, 0.0001392532, 8.552483e-05, 0, 0, 0,
  0, 0, 0, 5.851438e-09, 7.010658e-09, 7.010658e-09, 5.851438e-09, 0, 0, 0,
  0, 0, 1.763804e-08, 2.424815e-08, 2.875123e-08, 2.875123e-08, 2.424815e-08, 
    1.763804e-08, 0, 0,
  0, 1.763804e-08, 3.315868e-08, 2.900409e-08, 2.569869e-08, 2.569869e-08, 
    2.900409e-08, 3.315868e-08, 1.763804e-08, 0,
  5.851438e-09, 2.424815e-08, 2.900409e-08, 2.173926e-08, 1.616258e-08, 
    1.616258e-08, 2.173926e-08, 2.900409e-08, 2.424815e-08, 5.851438e-09,
  7.010658e-09, 2.875123e-08, 2.569869e-08, 1.616258e-08, 8.32039e-09, 
    8.32039e-09, 1.616258e-08, 2.569869e-08, 2.875123e-08, 7.010658e-09,
  7.010658e-09, 2.875123e-08, 2.569869e-08, 1.616258e-08, 8.32039e-09, 
    8.32039e-09, 1.616258e-08, 2.569869e-08, 2.875123e-08, 7.010658e-09,
  5.851438e-09, 2.424815e-08, 2.900409e-08, 2.173926e-08, 1.616258e-08, 
    1.616258e-08, 2.173926e-08, 2.900409e-08, 2.424815e-08, 5.851438e-09,
  0, 1.763804e-08, 3.315868e-08, 2.900409e-08, 2.569869e-08, 2.569869e-08, 
    2.900409e-08, 3.315868e-08, 1.763804e-08, 0,
  0, 0, 1.763804e-08, 2.424815e-08, 2.875123e-08, 2.875123e-08, 2.424815e-08, 
    1.763804e-08, 0, 0,
  0, 0, 0, 5.851438e-09, 7.010658e-09, 7.010658e-09, 5.851438e-09, 0, 0, 0,
  0, 0, 0, 0.0006154863, 0.0009428004, 0.0009428004, 0.0006154863, 0, 0, 0,
  0, 0, 0.0008176809, 0.002296266, 0.00352581, 0.00352581, 0.002296266, 
    0.0008176809, 0, 0,
  0, 0.0008176809, 0.0117573, 0.01075714, 0.009601971, 0.009601971, 
    0.01075714, 0.0117573, 0.0008176809, 0,
  0.0006154863, 0.002296266, 0.01075714, 0.006409943, 0.002547283, 
    0.002547283, 0.006409943, 0.01075714, 0.002296266, 0.0006154863,
  0.0009428004, 0.00352581, 0.009601971, 0.002547283, 0.0002127351, 
    0.0002127351, 0.002547283, 0.009601971, 0.00352581, 0.0009428004,
  0.0009428004, 0.00352581, 0.009601971, 0.002547283, 0.0002127351, 
    0.0002127351, 0.002547283, 0.009601971, 0.00352581, 0.0009428004,
  0.0006154863, 0.002296266, 0.01075714, 0.006409943, 0.002547283, 
    0.002547283, 0.006409943, 0.01075714, 0.002296266, 0.0006154863,
  0, 0.0008176809, 0.0117573, 0.01075714, 0.009601971, 0.009601971, 
    0.01075714, 0.0117573, 0.0008176809, 0,
  0, 0, 0.0008176809, 0.002296266, 0.00352581, 0.00352581, 0.002296266, 
    0.0008176809, 0, 0,
  0, 0, 0, 0.0006154863, 0.0009428004, 0.0009428004, 0.0006154863, 0, 0, 0,
  0, 0, 0, 0.0006027535, 0.0009313494, 0.0009313494, 0.0006027535, 0, 0, 0,
  0, 0, 0.000740111, 0.002248325, 0.0034784, 0.0034784, 0.002248325, 
    0.000740111, 0, 0,
  0, 0.000740111, 0.01165757, 0.01063941, 0.009475038, 0.009475038, 
    0.01063941, 0.01165757, 0.000740111, 0,
  0.0006027535, 0.002248325, 0.01063941, 0.006301843, 0.002466426, 
    0.002466426, 0.006301843, 0.01063941, 0.002248325, 0.0006027535,
  0.0009313494, 0.0034784, 0.009475038, 0.002466426, 0.0002003695, 
    0.0002003695, 0.002466426, 0.009475038, 0.0034784, 0.0009313494,
  0.0009313494, 0.0034784, 0.009475038, 0.002466426, 0.0002003695, 
    0.0002003695, 0.002466426, 0.009475038, 0.0034784, 0.0009313494,
  0.0006027535, 0.002248325, 0.01063941, 0.006301843, 0.002466426, 
    0.002466426, 0.006301843, 0.01063941, 0.002248325, 0.0006027535,
  0, 0.000740111, 0.01165757, 0.01063941, 0.009475038, 0.009475038, 
    0.01063941, 0.01165757, 0.000740111, 0,
  0, 0, 0.000740111, 0.002248325, 0.0034784, 0.0034784, 0.002248325, 
    0.000740111, 0, 0,
  0, 0, 0, 0.0006027535, 0.0009313494, 0.0009313494, 0.0006027535, 0, 0, 0,
  0, 0, 0, 0.0005701687, 0.000895333, 0.000895333, 0.0005701687, 0, 0, 0,
  0, 0, 0.0006008537, 0.002126917, 0.003341519, 0.003341519, 0.002126917, 
    0.0006008537, 0, 0,
  0, 0.0006008537, 0.01127949, 0.01027103, 0.009104954, 0.009104954, 
    0.01027103, 0.01127949, 0.0006008537, 0,
  0.0005701687, 0.002126917, 0.01027103, 0.005973883, 0.002264932, 
    0.002264932, 0.005973883, 0.01027103, 0.002126917, 0.0005701687,
  0.000895333, 0.003341519, 0.009104954, 0.002264932, 0.0001756543, 
    0.0001756543, 0.002264932, 0.009104954, 0.003341519, 0.000895333,
  0.000895333, 0.003341519, 0.009104954, 0.002264932, 0.0001756543, 
    0.0001756543, 0.002264932, 0.009104954, 0.003341519, 0.000895333,
  0.0005701687, 0.002126917, 0.01027103, 0.005973883, 0.002264932, 
    0.002264932, 0.005973883, 0.01027103, 0.002126917, 0.0005701687,
  0, 0.0006008537, 0.01127949, 0.01027103, 0.009104954, 0.009104954, 
    0.01027103, 0.01127949, 0.0006008537, 0,
  0, 0, 0.0006008537, 0.002126917, 0.003341519, 0.003341519, 0.002126917, 
    0.0006008537, 0, 0,
  0, 0, 0, 0.0005701687, 0.000895333, 0.000895333, 0.0005701687, 0, 0, 0,
  0, 0, 0, 0.0005161816, 0.000820153, 0.000820153, 0.0005161816, 0, 0, 0,
  0, 0, 0.000467052, 0.001925476, 0.003060083, 0.003060083, 0.001925476, 
    0.000467052, 0, 0,
  0, 0.000467052, 0.01042684, 0.009504506, 0.008408021, 0.008408021, 
    0.009504506, 0.01042684, 0.000467052, 0,
  0.0005161816, 0.001925476, 0.009504506, 0.005439742, 0.002002269, 
    0.002002269, 0.005439742, 0.009504506, 0.001925476, 0.0005161816,
  0.000820153, 0.003060083, 0.008408021, 0.002002269, 0.0001463965, 
    0.0001463965, 0.002002269, 0.008408021, 0.003060083, 0.000820153,
  0.000820153, 0.003060083, 0.008408021, 0.002002269, 0.0001463965, 
    0.0001463965, 0.002002269, 0.008408021, 0.003060083, 0.000820153,
  0.0005161816, 0.001925476, 0.009504506, 0.005439742, 0.002002269, 
    0.002002269, 0.005439742, 0.009504506, 0.001925476, 0.0005161816,
  0, 0.000467052, 0.01042684, 0.009504506, 0.008408021, 0.008408021, 
    0.009504506, 0.01042684, 0.000467052, 0,
  0, 0, 0.000467052, 0.001925476, 0.003060083, 0.003060083, 0.001925476, 
    0.000467052, 0, 0,
  0, 0, 0, 0.0005161816, 0.000820153, 0.000820153, 0.0005161816, 0, 0, 0,
  0, 0, 0, 0.0004432316, 0.0007097511, 0.0007097511, 0.0004432316, 0, 0, 0,
  0, 0, 0.0003507923, 0.001653381, 0.002647939, 0.002647939, 0.001653381, 
    0.0003507923, 0, 0,
  0, 0.0003507923, 0.009116829, 0.008327477, 0.007367987, 0.007367987, 
    0.008327477, 0.009116829, 0.0003507923, 0,
  0.0004432316, 0.001653381, 0.008327477, 0.004709304, 0.001698195, 
    0.001698195, 0.004709304, 0.008327477, 0.001653381, 0.0004432316,
  0.0007097511, 0.002647939, 0.007367987, 0.001698195, 0.00011795, 
    0.00011795, 0.001698195, 0.007367987, 0.002647939, 0.0007097511,
  0.0007097511, 0.002647939, 0.007367987, 0.001698195, 0.00011795, 
    0.00011795, 0.001698195, 0.007367987, 0.002647939, 0.0007097511,
  0.0004432316, 0.001653381, 0.008327477, 0.004709304, 0.001698195, 
    0.001698195, 0.004709304, 0.008327477, 0.001653381, 0.0004432316,
  0, 0.0003507923, 0.009116829, 0.008327477, 0.007367987, 0.007367987, 
    0.008327477, 0.009116829, 0.0003507923, 0,
  0, 0, 0.0003507923, 0.001653381, 0.002647939, 0.002647939, 0.001653381, 
    0.0003507923, 0, 0,
  0, 0, 0, 0.0004432316, 0.0007097511, 0.0007097511, 0.0004432316, 0, 0, 0,
  0, 0, 0, 0.000358204, 0.0005766553, 0.0005766553, 0.000358204, 0, 0, 0,
  0, 0, 0.0002528262, 0.001336272, 0.002151391, 0.002151391, 0.001336272, 
    0.0002528262, 0, 0,
  0, 0.0002528262, 0.00748521, 0.006850153, 0.006066464, 0.006066464, 
    0.006850153, 0.00748521, 0.0002528262, 0,
  0.000358204, 0.001336272, 0.006850153, 0.00383717, 0.001364885, 
    0.001364885, 0.00383717, 0.006850153, 0.001336272, 0.000358204,
  0.0005766553, 0.002151391, 0.006066464, 0.001364885, 9.177285e-05, 
    9.177285e-05, 0.001364885, 0.006066464, 0.002151391, 0.0005766553,
  0.0005766553, 0.002151391, 0.006066464, 0.001364885, 9.177285e-05, 
    9.177285e-05, 0.001364885, 0.006066464, 0.002151391, 0.0005766553,
  0.000358204, 0.001336272, 0.006850153, 0.00383717, 0.001364885, 
    0.001364885, 0.00383717, 0.006850153, 0.001336272, 0.000358204,
  0, 0.0002528262, 0.00748521, 0.006850153, 0.006066464, 0.006066464, 
    0.006850153, 0.00748521, 0.0002528262, 0,
  0, 0, 0.0002528262, 0.001336272, 0.002151391, 0.002151391, 0.001336272, 
    0.0002528262, 0, 0,
  0, 0, 0, 0.000358204, 0.0005766553, 0.0005766553, 0.000358204, 0, 0, 0,
  0, 0, 0, 0.00026761, 0.0004323024, 0.0004323024, 0.00026761, 0, 0, 0,
  0, 0, 0.0001719894, 0.000998384, 0.001612911, 0.001612911, 0.000998384, 
    0.0001719894, 0, 0,
  0, 0.0001719894, 0.005671083, 0.005197524, 0.004607539, 0.004607539, 
    0.005197524, 0.005671083, 0.0001719894, 0,
  0.00026761, 0.000998384, 0.005197524, 0.002887747, 0.001017328, 
    0.001017328, 0.002887747, 0.005197524, 0.000998384, 0.00026761,
  0.0004323024, 0.001612911, 0.004607539, 0.001017328, 6.728976e-05, 
    6.728976e-05, 0.001017328, 0.004607539, 0.001612911, 0.0004323024,
  0.0004323024, 0.001612911, 0.004607539, 0.001017328, 6.728976e-05, 
    6.728976e-05, 0.001017328, 0.004607539, 0.001612911, 0.0004323024,
  0.00026761, 0.000998384, 0.005197524, 0.002887747, 0.001017328, 
    0.001017328, 0.002887747, 0.005197524, 0.000998384, 0.00026761,
  0, 0.0001719894, 0.005671083, 0.005197524, 0.004607539, 0.004607539, 
    0.005197524, 0.005671083, 0.0001719894, 0,
  0, 0, 0.0001719894, 0.000998384, 0.001612911, 0.001612911, 0.000998384, 
    0.0001719894, 0, 0,
  0, 0, 0, 0.00026761, 0.0004323024, 0.0004323024, 0.00026761, 0, 0, 0,
  0, 0, 0, 0.0001760609, 0.0002850214, 0.0002850214, 0.0001760609, 0, 0, 0,
  0, 0, 0.0001049547, 0.0006568938, 0.001063483, 0.001063483, 0.0006568938, 
    0.0001049547, 0, 0,
  0, 0.0001049547, 0.003780114, 0.003469298, 0.003078709, 0.003078709, 
    0.003469298, 0.003780114, 0.0001049547, 0,
  0.0001760609, 0.0006568938, 0.003469298, 0.001913728, 0.0006691327, 
    0.0006691327, 0.001913728, 0.003469298, 0.0006568938, 0.0001760609,
  0.0002850214, 0.001063483, 0.003078709, 0.0006691327, 4.400047e-05, 
    4.400047e-05, 0.0006691327, 0.003078709, 0.001063483, 0.0002850214,
  0.0002850214, 0.001063483, 0.003078709, 0.0006691327, 4.400047e-05, 
    4.400047e-05, 0.0006691327, 0.003078709, 0.001063483, 0.0002850214,
  0.0001760609, 0.0006568938, 0.003469298, 0.001913728, 0.0006691327, 
    0.0006691327, 0.001913728, 0.003469298, 0.0006568938, 0.0001760609,
  0, 0.0001049547, 0.003780114, 0.003469298, 0.003078709, 0.003078709, 
    0.003469298, 0.003780114, 0.0001049547, 0,
  0, 0, 0.0001049547, 0.0006568938, 0.001063483, 0.001063483, 0.0006568938, 
    0.0001049547, 0, 0,
  0, 0, 0, 0.0001760609, 0.0002850214, 0.0002850214, 0.0001760609, 0, 0, 0,
  0, 0, 0, 8.63148e-05, 0.000140021, 0.000140021, 8.63148e-05, 0, 0, 0,
  0, 0, 4.803922e-05, 0.000322081, 0.0005225019, 0.0005225019, 0.000322081, 
    4.803922e-05, 0, 0,
  0, 4.803922e-05, 0.001878512, 0.00172877, 0.001537071, 0.001537071, 
    0.00172877, 0.001878512, 4.803922e-05, 0,
  8.63148e-05, 0.000322081, 0.00172877, 0.0009491512, 0.0003296222, 
    0.0003296222, 0.0009491512, 0.00172877, 0.000322081, 8.63148e-05,
  0.000140021, 0.0005225019, 0.001537071, 0.0003296222, 2.168196e-05, 
    2.168196e-05, 0.0003296222, 0.001537071, 0.0005225019, 0.000140021,
  0.000140021, 0.0005225019, 0.001537071, 0.0003296222, 2.168196e-05, 
    2.168196e-05, 0.0003296222, 0.001537071, 0.0005225019, 0.000140021,
  8.63148e-05, 0.000322081, 0.00172877, 0.0009491512, 0.0003296222, 
    0.0003296222, 0.0009491512, 0.00172877, 0.000322081, 8.63148e-05,
  0, 4.803922e-05, 0.001878512, 0.00172877, 0.001537071, 0.001537071, 
    0.00172877, 0.001878512, 4.803922e-05, 0,
  0, 0, 4.803922e-05, 0.000322081, 0.0005225019, 0.0005225019, 0.000322081, 
    4.803922e-05, 0, 0,
  0, 0, 0, 8.63148e-05, 0.000140021, 0.000140021, 8.63148e-05, 0, 0, 0,
  0, 0, 0, 5.854663e-09, 7.011049e-09, 7.011049e-09, 5.854663e-09, 0, 0, 0,
  0, 0, 1.766774e-08, 2.427772e-08, 2.877424e-08, 2.877424e-08, 2.427772e-08, 
    1.766774e-08, 0, 0,
  0, 1.766774e-08, 3.314915e-08, 2.895513e-08, 2.562989e-08, 2.562989e-08, 
    2.895513e-08, 3.314915e-08, 1.766774e-08, 0,
  5.854663e-09, 2.427772e-08, 2.895513e-08, 2.17148e-08, 1.616976e-08, 
    1.616976e-08, 2.17148e-08, 2.895513e-08, 2.427772e-08, 5.854663e-09,
  7.011049e-09, 2.877424e-08, 2.562989e-08, 1.616976e-08, 8.349289e-09, 
    8.349289e-09, 1.616976e-08, 2.562989e-08, 2.877424e-08, 7.011049e-09,
  7.011049e-09, 2.877424e-08, 2.562989e-08, 1.616976e-08, 8.349289e-09, 
    8.349289e-09, 1.616976e-08, 2.562989e-08, 2.877424e-08, 7.011049e-09,
  5.854663e-09, 2.427772e-08, 2.895513e-08, 2.17148e-08, 1.616976e-08, 
    1.616976e-08, 2.17148e-08, 2.895513e-08, 2.427772e-08, 5.854663e-09,
  0, 1.766774e-08, 3.314915e-08, 2.895513e-08, 2.562989e-08, 2.562989e-08, 
    2.895513e-08, 3.314915e-08, 1.766774e-08, 0,
  0, 0, 1.766774e-08, 2.427772e-08, 2.877424e-08, 2.877424e-08, 2.427772e-08, 
    1.766774e-08, 0, 0,
  0, 0, 0, 5.854663e-09, 7.011049e-09, 7.011049e-09, 5.854663e-09, 0, 0, 0,
  0, 0, 0, 0.0005094535, 0.0009715963, 0.0009715963, 0.0005094535, 0, 0, 0,
  0, 0.0001738648, 0.0007657561, 0.001901258, 0.003633362, 0.003633362, 
    0.001901258, 0.0007657561, 0.0001738648, 0,
  0, 0.0007657561, 0.003310008, 0.01048081, 0.009588317, 0.009588317, 
    0.01048081, 0.003310008, 0.0007657561, 0,
  0.0005094535, 0.001901258, 0.01048081, 0.006015534, 0.002596516, 
    0.002596516, 0.006015534, 0.01048081, 0.001901258, 0.0005094535,
  0.0009715963, 0.003633362, 0.009588317, 0.002596516, 0.0002088121, 
    0.0002088121, 0.002596516, 0.009588317, 0.003633362, 0.0009715963,
  0.0009715963, 0.003633362, 0.009588317, 0.002596516, 0.0002088121, 
    0.0002088121, 0.002596516, 0.009588317, 0.003633362, 0.0009715963,
  0.0005094535, 0.001901258, 0.01048081, 0.006015534, 0.002596516, 
    0.002596516, 0.006015534, 0.01048081, 0.001901258, 0.0005094535,
  0, 0.0007657561, 0.003310008, 0.01048081, 0.009588317, 0.009588317, 
    0.01048081, 0.003310008, 0.0007657561, 0,
  0, 0.0001738648, 0.0007657561, 0.001901258, 0.003633362, 0.003633362, 
    0.001901258, 0.0007657561, 0.0001738648, 0,
  0, 0, 0, 0.0005094535, 0.0009715963, 0.0009715963, 0.0005094535, 0, 0, 0,
  0, 0, 0, 0.000495396, 0.0009604159, 0.0009604159, 0.000495396, 0, 0, 0,
  0, 0.0001770358, 0.0007632556, 0.001849997, 0.003586487, 0.003586487, 
    0.001849997, 0.0007632556, 0.0001770358, 0,
  0, 0.0007632556, 0.003246959, 0.01036223, 0.009462952, 0.009462952, 
    0.01036223, 0.003246959, 0.0007632556, 0,
  0.000495396, 0.001849997, 0.01036223, 0.005932671, 0.002511997, 
    0.002511997, 0.005932671, 0.01036223, 0.001849997, 0.000495396,
  0.0009604159, 0.003586487, 0.009462952, 0.002511997, 0.0001970624, 
    0.0001970624, 0.002511997, 0.009462952, 0.003586487, 0.0009604159,
  0.0009604159, 0.003586487, 0.009462952, 0.002511997, 0.0001970624, 
    0.0001970624, 0.002511997, 0.009462952, 0.003586487, 0.0009604159,
  0.000495396, 0.001849997, 0.01036223, 0.005932671, 0.002511997, 
    0.002511997, 0.005932671, 0.01036223, 0.001849997, 0.000495396,
  0, 0.0007632556, 0.003246959, 0.01036223, 0.009462952, 0.009462952, 
    0.01036223, 0.003246959, 0.0007632556, 0,
  0, 0.0001770358, 0.0007632556, 0.001849997, 0.003586487, 0.003586487, 
    0.001849997, 0.0007632556, 0.0001770358, 0,
  0, 0, 0, 0.000495396, 0.0009604159, 0.0009604159, 0.000495396, 0, 0, 0,
  0, 0, 0, 0.0004624494, 0.00092431, 0.00092431, 0.0004624494, 0, 0, 0,
  0, 0.0001765596, 0.0007412257, 0.001727641, 0.003449111, 0.003449111, 
    0.001727641, 0.0007412257, 0.0001765596, 0,
  0, 0.0007412257, 0.003088127, 0.009997355, 0.009096014, 0.009096014, 
    0.009997355, 0.003088127, 0.0007412257, 0,
  0.0004624494, 0.001727641, 0.009997355, 0.005652009, 0.002305039, 
    0.002305039, 0.005652009, 0.009997355, 0.001727641, 0.0004624494,
  0.00092431, 0.003449111, 0.009096014, 0.002305039, 0.0001729962, 
    0.0001729962, 0.002305039, 0.009096014, 0.003449111, 0.00092431,
  0.00092431, 0.003449111, 0.009096014, 0.002305039, 0.0001729962, 
    0.0001729962, 0.002305039, 0.009096014, 0.003449111, 0.00092431,
  0.0004624494, 0.001727641, 0.009997355, 0.005652009, 0.002305039, 
    0.002305039, 0.005652009, 0.009997355, 0.001727641, 0.0004624494,
  0, 0.0007412257, 0.003088127, 0.009997355, 0.009096014, 0.009096014, 
    0.009997355, 0.003088127, 0.0007412257, 0,
  0, 0.0001765596, 0.0007412257, 0.001727641, 0.003449111, 0.003449111, 
    0.001727641, 0.0007412257, 0.0001765596, 0,
  0, 0, 0, 0.0004624494, 0.00092431, 0.00092431, 0.0004624494, 0, 0, 0,
  0, 0, 0, 0.000414066, 0.0008475719, 0.0008475719, 0.000414066, 0, 0, 0,
  0, 0.000166133, 0.0006850364, 0.001546742, 0.003161913, 0.003161913, 
    0.001546742, 0.0006850364, 0.000166133, 0,
  0, 0.0006850364, 0.0028119, 0.009253463, 0.008401131, 0.008401131, 
    0.009253463, 0.0028119, 0.0006850364, 0,
  0.000414066, 0.001546742, 0.009253463, 0.005167077, 0.002037211, 
    0.002037211, 0.005167077, 0.009253463, 0.001546742, 0.000414066,
  0.0008475719, 0.003161913, 0.008401131, 0.002037211, 0.0001441602, 
    0.0001441602, 0.002037211, 0.008401131, 0.003161913, 0.0008475719,
  0.0008475719, 0.003161913, 0.008401131, 0.002037211, 0.0001441602, 
    0.0001441602, 0.002037211, 0.008401131, 0.003161913, 0.0008475719,
  0.000414066, 0.001546742, 0.009253463, 0.005167077, 0.002037211, 
    0.002037211, 0.005167077, 0.009253463, 0.001546742, 0.000414066,
  0, 0.0006850364, 0.0028119, 0.009253463, 0.008401131, 0.008401131, 
    0.009253463, 0.0028119, 0.0006850364, 0,
  0, 0.000166133, 0.0006850364, 0.001546742, 0.003161913, 0.003161913, 
    0.001546742, 0.0006850364, 0.000166133, 0,
  0, 0, 0, 0.000414066, 0.0008475719, 0.0008475719, 0.000414066, 0, 0, 0,
  0, 0, 0, 0.0003528663, 0.0007340594, 0.0007340594, 0.0003528663, 0, 0, 0,
  0, 0.0001464571, 0.0005971373, 0.001317893, 0.002738278, 0.002738278, 
    0.001317893, 0.0005971373, 0.0001464571, 0,
  0, 0.0005971373, 0.00242749, 0.008114112, 0.00736268, 0.00736268, 
    0.008114112, 0.00242749, 0.0005971373, 0,
  0.0003528663, 0.001317893, 0.008114112, 0.00448683, 0.001727467, 
    0.001727467, 0.00448683, 0.008114112, 0.001317893, 0.0003528663,
  0.0007340594, 0.002738278, 0.00736268, 0.001727467, 0.0001161502, 
    0.0001161502, 0.001727467, 0.00736268, 0.002738278, 0.0007340594,
  0.0007340594, 0.002738278, 0.00736268, 0.001727467, 0.0001161502, 
    0.0001161502, 0.001727467, 0.00736268, 0.002738278, 0.0007340594,
  0.0003528663, 0.001317893, 0.008114112, 0.00448683, 0.001727467, 
    0.001727467, 0.00448683, 0.008114112, 0.001317893, 0.0003528663,
  0, 0.0005971373, 0.00242749, 0.008114112, 0.00736268, 0.00736268, 
    0.008114112, 0.00242749, 0.0005971373, 0,
  0, 0.0001464571, 0.0005971373, 0.001317893, 0.002738278, 0.002738278, 
    0.001317893, 0.0005971373, 0.0001464571, 0,
  0, 0, 0, 0.0003528663, 0.0007340594, 0.0007340594, 0.0003528663, 0, 0, 0,
  0, 0, 0, 0.0002836539, 0.0005967911, 0.0005967911, 0.0002836539, 0, 0, 0,
  0, 0.0001206066, 0.0004881136, 0.001059214, 0.002226282, 0.002226282, 
    0.001059214, 0.0004881136, 0.0001206066, 0,
  0, 0.0004881136, 0.001971457, 0.006681798, 0.00606292, 0.00606292, 
    0.006681798, 0.001971457, 0.0004881136, 0,
  0.0002836539, 0.001059214, 0.006681798, 0.003664744, 0.001388144, 
    0.001388144, 0.003664744, 0.006681798, 0.001059214, 0.0002836539,
  0.0005967911, 0.002226282, 0.00606292, 0.001388144, 9.042394e-05, 
    9.042394e-05, 0.001388144, 0.00606292, 0.002226282, 0.0005967911,
  0.0005967911, 0.002226282, 0.00606292, 0.001388144, 9.042394e-05, 
    9.042394e-05, 0.001388144, 0.00606292, 0.002226282, 0.0005967911,
  0.0002836539, 0.001059214, 0.006681798, 0.003664744, 0.001388144, 
    0.001388144, 0.003664744, 0.006681798, 0.001059214, 0.0002836539,
  0, 0.0004881136, 0.001971457, 0.006681798, 0.00606292, 0.00606292, 
    0.006681798, 0.001971457, 0.0004881136, 0,
  0, 0.0001206066, 0.0004881136, 0.001059214, 0.002226282, 0.002226282, 
    0.001059214, 0.0004881136, 0.0001206066, 0,
  0, 0, 0, 0.0002836539, 0.0005967911, 0.0005967911, 0.0002836539, 0, 0, 0,
  0, 0, 0, 0.0002110996, 0.0004476599, 0.0004476599, 0.0002110996, 0, 0, 0,
  0, 9.134485e-05, 0.0003678787, 0.0007881612, 0.001670075, 0.001670075, 
    0.0007881612, 0.0003678787, 9.134485e-05, 0,
  0, 0.0003678787, 0.001479404, 0.005076186, 0.004606068, 0.004606068, 
    0.005076186, 0.001479404, 0.0003678787, 0,
  0.0002110996, 0.0007881612, 0.005076186, 0.002763638, 0.001034584, 
    0.001034584, 0.002763638, 0.005076186, 0.0007881612, 0.0002110996,
  0.0004476599, 0.001670075, 0.004606068, 0.001034584, 6.636605e-05, 
    6.636605e-05, 0.001034584, 0.004606068, 0.001670075, 0.0004476599,
  0.0004476599, 0.001670075, 0.004606068, 0.001034584, 6.636605e-05, 
    6.636605e-05, 0.001034584, 0.004606068, 0.001670075, 0.0004476599,
  0.0002110996, 0.0007881612, 0.005076186, 0.002763638, 0.001034584, 
    0.001034584, 0.002763638, 0.005076186, 0.0007881612, 0.0002110996,
  0, 0.0003678787, 0.001479404, 0.005076186, 0.004606068, 0.004606068, 
    0.005076186, 0.001479404, 0.0003678787, 0,
  0, 9.134485e-05, 0.0003678787, 0.0007881612, 0.001670075, 0.001670075, 
    0.0007881612, 0.0003678787, 9.134485e-05, 0,
  0, 0, 0, 0.0002110996, 0.0004476599, 0.0004476599, 0.0002110996, 0, 0, 0,
  0, 0, 0, 0.0001384695, 0.0002953201, 0.0002953201, 0.0001384695, 0, 0, 0,
  0, 6.070226e-05, 0.0002436762, 0.0005169166, 0.001101846, 0.001101846, 
    0.0005169166, 0.0002436762, 6.070226e-05, 0,
  0, 0.0002436762, 0.0009771216, 0.003393139, 0.003079294, 0.003079294, 
    0.003393139, 0.0009771216, 0.0002436762, 0,
  0.0001384695, 0.0005169166, 0.003393139, 0.001835072, 0.0006806147, 
    0.0006806147, 0.001835072, 0.003393139, 0.0005169166, 0.0001384695,
  0.0002953201, 0.001101846, 0.003079294, 0.0006806147, 4.345326e-05, 
    4.345326e-05, 0.0006806147, 0.003079294, 0.001101846, 0.0002953201,
  0.0002953201, 0.001101846, 0.003079294, 0.0006806147, 4.345326e-05, 
    4.345326e-05, 0.0006806147, 0.003079294, 0.001101846, 0.0002953201,
  0.0001384695, 0.0005169166, 0.003393139, 0.001835072, 0.0006806147, 
    0.0006806147, 0.001835072, 0.003393139, 0.0005169166, 0.0001384695,
  0, 0.0002436762, 0.0009771216, 0.003393139, 0.003079294, 0.003079294, 
    0.003393139, 0.0009771216, 0.0002436762, 0,
  0, 6.070226e-05, 0.0002436762, 0.0005169166, 0.001101846, 0.001101846, 
    0.0005169166, 0.0002436762, 6.070226e-05, 0,
  0, 0, 0, 0.0001384695, 0.0002953201, 0.0002953201, 0.0001384695, 0, 0, 0,
  0, 0, 0, 6.768364e-05, 0.0001451609, 0.0001451609, 6.768364e-05, 0, 0, 0,
  0, 2.99955e-05, 0.0001201263, 0.000252635, 0.0005416647, 0.0005416647, 
    0.000252635, 0.0001201263, 2.99955e-05, 0,
  0, 0.0001201263, 0.0004807284, 0.0016931, 0.001538518, 0.001538518, 
    0.0016931, 0.0004807284, 0.0001201263, 0,
  6.768364e-05, 0.000252635, 0.0016931, 0.0009120474, 0.0003355041, 
    0.0003355041, 0.0009120474, 0.0016931, 0.000252635, 6.768364e-05,
  0.0001451609, 0.0005416647, 0.001538518, 0.0003355041, 2.14452e-05, 
    2.14452e-05, 0.0003355041, 0.001538518, 0.0005416647, 0.0001451609,
  0.0001451609, 0.0005416647, 0.001538518, 0.0003355041, 2.14452e-05, 
    2.14452e-05, 0.0003355041, 0.001538518, 0.0005416647, 0.0001451609,
  6.768364e-05, 0.000252635, 0.0016931, 0.0009120474, 0.0003355041, 
    0.0003355041, 0.0009120474, 0.0016931, 0.000252635, 6.768364e-05,
  0, 0.0001201263, 0.0004807284, 0.0016931, 0.001538518, 0.001538518, 
    0.0016931, 0.0004807284, 0.0001201263, 0,
  0, 2.99955e-05, 0.0001201263, 0.000252635, 0.0005416647, 0.0005416647, 
    0.000252635, 0.0001201263, 2.99955e-05, 0,
  0, 0, 0, 6.768364e-05, 0.0001451609, 0.0001451609, 6.768364e-05, 0, 0, 0,
  0, 0, 0, 5.872243e-09, 7.011028e-09, 7.011028e-09, 5.872243e-09, 0, 0, 0,
  0, 3.280666e-09, 6.249122e-09, 2.431012e-08, 2.880439e-08, 2.880439e-08, 
    2.431012e-08, 6.249122e-09, 3.280666e-09, 0,
  0, 6.249122e-09, 2.657537e-08, 2.879584e-08, 2.555656e-08, 2.555656e-08, 
    2.879584e-08, 2.657537e-08, 6.249122e-09, 0,
  5.872243e-09, 2.431012e-08, 2.879584e-08, 2.135364e-08, 1.622879e-08, 
    1.622879e-08, 2.135364e-08, 2.879584e-08, 2.431012e-08, 5.872243e-09,
  7.011028e-09, 2.880439e-08, 2.555656e-08, 1.622879e-08, 8.358248e-09, 
    8.358248e-09, 1.622879e-08, 2.555656e-08, 2.880439e-08, 7.011028e-09,
  7.011028e-09, 2.880439e-08, 2.555656e-08, 1.622879e-08, 8.358248e-09, 
    8.358248e-09, 1.622879e-08, 2.555656e-08, 2.880439e-08, 7.011028e-09,
  5.872243e-09, 2.431012e-08, 2.879584e-08, 2.135364e-08, 1.622879e-08, 
    1.622879e-08, 2.135364e-08, 2.879584e-08, 2.431012e-08, 5.872243e-09,
  0, 6.249122e-09, 2.657537e-08, 2.879584e-08, 2.555656e-08, 2.555656e-08, 
    2.879584e-08, 2.657537e-08, 6.249122e-09, 0,
  0, 3.280666e-09, 6.249122e-09, 2.431012e-08, 2.880439e-08, 2.880439e-08, 
    2.431012e-08, 6.249122e-09, 3.280666e-09, 0,
  0, 0, 0, 5.872243e-09, 7.011028e-09, 7.011028e-09, 5.872243e-09, 0, 0, 0,
  0, 0, 0, 0.0005135111, 0.000975395, 0.000975395, 0.0005135111, 0, 0, 0,
  0, 0.0001742384, 0.0007684355, 0.001916463, 0.003647718, 0.003647718, 
    0.001916463, 0.0007684355, 0.0001742384, 0,
  0, 0.0007684355, 0.003324748, 0.01045375, 0.009532276, 0.009532276, 
    0.01045375, 0.003324748, 0.0007684355, 0,
  0.0005135111, 0.001916463, 0.01045375, 0.00598867, 0.002600763, 
    0.002600763, 0.00598867, 0.01045375, 0.001916463, 0.0005135111,
  0.000975395, 0.003647718, 0.009532276, 0.002600763, 0.0002123007, 
    0.0002123007, 0.002600763, 0.009532276, 0.003647718, 0.000975395,
  0.000975395, 0.003647718, 0.009532276, 0.002600763, 0.0002123007, 
    0.0002123007, 0.002600763, 0.009532276, 0.003647718, 0.000975395,
  0.0005135111, 0.001916463, 0.01045375, 0.00598867, 0.002600763, 
    0.002600763, 0.00598867, 0.01045375, 0.001916463, 0.0005135111,
  0, 0.0007684355, 0.003324748, 0.01045375, 0.009532276, 0.009532276, 
    0.01045375, 0.003324748, 0.0007684355, 0,
  0, 0.0001742384, 0.0007684355, 0.001916463, 0.003647718, 0.003647718, 
    0.001916463, 0.0007684355, 0.0001742384, 0,
  0, 0, 0, 0.0005135111, 0.000975395, 0.000975395, 0.0005135111, 0, 0, 0,
  0, 0, 0, 0.0004994313, 0.0009642431, 0.0009642431, 0.0004994313, 0, 0, 0,
  0, 0.000177459, 0.0007660275, 0.001865088, 0.003600866, 0.003600866, 
    0.001865088, 0.0007660275, 0.000177459, 0,
  0, 0.0007660275, 0.003261694, 0.01033576, 0.009408205, 0.009408205, 
    0.01033576, 0.003261694, 0.0007660275, 0,
  0.0004994313, 0.001865088, 0.01033576, 0.005906021, 0.002516394, 
    0.002516394, 0.005906021, 0.01033576, 0.001865088, 0.0004994313,
  0.0009642431, 0.003600866, 0.009408205, 0.002516394, 0.000200392, 
    0.000200392, 0.002516394, 0.009408205, 0.003600866, 0.0009642431,
  0.0009642431, 0.003600866, 0.009408205, 0.002516394, 0.000200392, 
    0.000200392, 0.002516394, 0.009408205, 0.003600866, 0.0009642431,
  0.0004994313, 0.001865088, 0.01033576, 0.005906021, 0.002516394, 
    0.002516394, 0.005906021, 0.01033576, 0.001865088, 0.0004994313,
  0, 0.0007660275, 0.003261694, 0.01033576, 0.009408205, 0.009408205, 
    0.01033576, 0.003261694, 0.0007660275, 0,
  0, 0.000177459, 0.0007660275, 0.001865088, 0.003600866, 0.003600866, 
    0.001865088, 0.0007660275, 0.000177459, 0,
  0, 0, 0, 0.0004994313, 0.0009642431, 0.0009642431, 0.0004994313, 0, 0, 0,
  0, 0, 0, 0.0004663947, 0.0009280923, 0.0009280923, 0.0004663947, 0, 0, 0,
  0, 0.000177049, 0.0007440911, 0.001742378, 0.003463273, 0.003463273, 
    0.001742378, 0.0007440911, 0.000177049, 0,
  0, 0.0007440911, 0.003102627, 0.009972387, 0.009044145, 0.009044145, 
    0.009972387, 0.003102627, 0.0007440911, 0,
  0.0004663947, 0.001742378, 0.009972387, 0.005626449, 0.002309881, 
    0.002309881, 0.005626449, 0.009972387, 0.001742378, 0.0004663947,
  0.0009280923, 0.003463273, 0.009044145, 0.002309881, 0.0001759276, 
    0.0001759276, 0.002309881, 0.009044145, 0.003463273, 0.0009280923,
  0.0009280923, 0.003463273, 0.009044145, 0.002309881, 0.0001759276, 
    0.0001759276, 0.002309881, 0.009044145, 0.003463273, 0.0009280923,
  0.0004663947, 0.001742378, 0.009972387, 0.005626449, 0.002309881, 
    0.002309881, 0.005626449, 0.009972387, 0.001742378, 0.0004663947,
  0, 0.0007440911, 0.003102627, 0.009972387, 0.009044145, 0.009044145, 
    0.009972387, 0.003102627, 0.0007440911, 0,
  0, 0.000177049, 0.0007440911, 0.001742378, 0.003463273, 0.003463273, 
    0.001742378, 0.0007440911, 0.000177049, 0,
  0, 0, 0, 0.0004663947, 0.0009280923, 0.0009280923, 0.0004663947, 0, 0, 0,
  0, 0, 0, 0.0004177446, 0.0008511285, 0.0008511285, 0.0004177446, 0, 0, 0,
  0, 0.0001666484, 0.000687848, 0.001560473, 0.00317521, 0.00317521, 
    0.001560473, 0.000687848, 0.0001666484, 0,
  0, 0.000687848, 0.00282562, 0.009231299, 0.008353945, 0.008353945, 
    0.009231299, 0.00282562, 0.000687848, 0,
  0.0004177446, 0.001560473, 0.009231299, 0.005143668, 0.002042309, 
    0.002042309, 0.005143668, 0.009231299, 0.001560473, 0.0004177446,
  0.0008511285, 0.00317521, 0.008353945, 0.002042309, 0.0001466312, 
    0.0001466312, 0.002042309, 0.008353945, 0.00317521, 0.0008511285,
  0.0008511285, 0.00317521, 0.008353945, 0.002042309, 0.0001466312, 
    0.0001466312, 0.002042309, 0.008353945, 0.00317521, 0.0008511285,
  0.0004177446, 0.001560473, 0.009231299, 0.005143668, 0.002042309, 
    0.002042309, 0.005143668, 0.009231299, 0.001560473, 0.0004177446,
  0, 0.000687848, 0.00282562, 0.009231299, 0.008353945, 0.008353945, 
    0.009231299, 0.00282562, 0.000687848, 0,
  0, 0.0001666484, 0.000687848, 0.001560473, 0.00317521, 0.00317521, 
    0.001560473, 0.000687848, 0.0001666484, 0,
  0, 0, 0, 0.0004177446, 0.0008511285, 0.0008511285, 0.0004177446, 0, 0, 0,
  0, 0, 0, 0.0003561142, 0.0007372297, 0.0007372297, 0.0003561142, 0, 0, 0,
  0, 0.000146956, 0.000599739, 0.001330014, 0.002750121, 0.002750121, 
    0.001330014, 0.000599739, 0.000146956, 0,
  0, 0.000599739, 0.002439864, 0.008096056, 0.007322218, 0.007322218, 
    0.008096056, 0.002439864, 0.000599739, 0,
  0.0003561142, 0.001330014, 0.008096056, 0.004466613, 0.001732403, 
    0.001732403, 0.004466613, 0.008096056, 0.001330014, 0.0003561142,
  0.0007372297, 0.002750121, 0.007322218, 0.001732403, 0.0001181813, 
    0.0001181813, 0.001732403, 0.007322218, 0.002750121, 0.0007372297,
  0.0007372297, 0.002750121, 0.007322218, 0.001732403, 0.0001181813, 
    0.0001181813, 0.001732403, 0.007322218, 0.002750121, 0.0007372297,
  0.0003561142, 0.001330014, 0.008096056, 0.004466613, 0.001732403, 
    0.001732403, 0.004466613, 0.008096056, 0.001330014, 0.0003561142,
  0, 0.000599739, 0.002439864, 0.008096056, 0.007322218, 0.007322218, 
    0.008096056, 0.002439864, 0.000599739, 0,
  0, 0.000146956, 0.000599739, 0.001330014, 0.002750121, 0.002750121, 
    0.001330014, 0.000599739, 0.000146956, 0,
  0, 0, 0, 0.0003561142, 0.0007372297, 0.0007372297, 0.0003561142, 0, 0, 0,
  0, 0, 0, 0.0002863611, 0.0005994588, 0.0005994588, 0.0002863611, 0, 0, 0,
  0, 0.0001210555, 0.0004903803, 0.001069315, 0.002236242, 0.002236242, 
    0.001069315, 0.0004903803, 0.0001210555, 0,
  0, 0.0004903803, 0.001982026, 0.006668716, 0.006030808, 0.006030808, 
    0.006668716, 0.001982026, 0.0004903803, 0,
  0.0002863611, 0.001069315, 0.006668716, 0.003648539, 0.001392569, 
    0.001392569, 0.003648539, 0.006668716, 0.001069315, 0.0002863611,
  0.0005994588, 0.002236242, 0.006030808, 0.001392569, 9.203804e-05, 
    9.203804e-05, 0.001392569, 0.006030808, 0.002236242, 0.0005994588,
  0.0005994588, 0.002236242, 0.006030808, 0.001392569, 9.203804e-05, 
    9.203804e-05, 0.001392569, 0.006030808, 0.002236242, 0.0005994588,
  0.0002863611, 0.001069315, 0.006668716, 0.003648539, 0.001392569, 
    0.001392569, 0.003648539, 0.006668716, 0.001069315, 0.0002863611,
  0, 0.0004903803, 0.001982026, 0.006668716, 0.006030808, 0.006030808, 
    0.006668716, 0.001982026, 0.0004903803, 0,
  0, 0.0001210555, 0.0004903803, 0.001069315, 0.002236242, 0.002236242, 
    0.001069315, 0.0004903803, 0.0001210555, 0,
  0, 0, 0, 0.0002863611, 0.0005994588, 0.0005994588, 0.0002863611, 0, 0, 0,
  0, 0, 0, 0.0002131898, 0.0004497514, 0.0004497514, 0.0002131898, 0, 0, 0,
  0, 9.171638e-05, 0.0003697058, 0.0007959589, 0.001677881, 0.001677881, 
    0.0007959589, 0.0003697058, 9.171638e-05, 0,
  0, 0.0003697058, 0.001487781, 0.005068295, 0.004583258, 0.004583258, 
    0.005068295, 0.001487781, 0.0003697058, 0,
  0.0002131898, 0.0007959589, 0.005068295, 0.002752012, 0.001038272, 
    0.001038272, 0.002752012, 0.005068295, 0.0007959589, 0.0002131898,
  0.0004497514, 0.001677881, 0.004583258, 0.001038272, 6.75785e-05, 
    6.75785e-05, 0.001038272, 0.004583258, 0.001677881, 0.0004497514,
  0.0004497514, 0.001677881, 0.004583258, 0.001038272, 6.75785e-05, 
    6.75785e-05, 0.001038272, 0.004583258, 0.001677881, 0.0004497514,
  0.0002131898, 0.0007959589, 0.005068295, 0.002752012, 0.001038272, 
    0.001038272, 0.002752012, 0.005068295, 0.0007959589, 0.0002131898,
  0, 0.0003697058, 0.001487781, 0.005068295, 0.004583258, 0.004583258, 
    0.005068295, 0.001487781, 0.0003697058, 0,
  0, 9.171638e-05, 0.0003697058, 0.0007959589, 0.001677881, 0.001677881, 
    0.0007959589, 0.0003697058, 9.171638e-05, 0,
  0, 0, 0, 0.0002131898, 0.0004497514, 0.0004497514, 0.0002131898, 0, 0, 0,
  0, 0, 0, 0.0001398786, 0.0002967776, 0.0002967776, 0.0001398786, 0, 0, 0,
  0, 6.097033e-05, 0.0002449627, 0.0005221736, 0.001107285, 0.001107285, 
    0.0005221736, 0.0002449627, 6.097033e-05, 0,
  0, 0.0002449627, 0.0009829302, 0.003389748, 0.003065823, 0.003065823, 
    0.003389748, 0.0009829302, 0.0002449627, 0,
  0.0001398786, 0.0005221736, 0.003389748, 0.001828278, 0.0006834217, 
    0.0006834217, 0.001828278, 0.003389748, 0.0005221736, 0.0001398786,
  0.0002967776, 0.001107285, 0.003065823, 0.0006834217, 4.427295e-05, 
    4.427295e-05, 0.0006834217, 0.003065823, 0.001107285, 0.0002967776,
  0.0002967776, 0.001107285, 0.003065823, 0.0006834217, 4.427295e-05, 
    4.427295e-05, 0.0006834217, 0.003065823, 0.001107285, 0.0002967776,
  0.0001398786, 0.0005221736, 0.003389748, 0.001828278, 0.0006834217, 
    0.0006834217, 0.001828278, 0.003389748, 0.0005221736, 0.0001398786,
  0, 0.0002449627, 0.0009829302, 0.003389748, 0.003065823, 0.003065823, 
    0.003389748, 0.0009829302, 0.0002449627, 0,
  0, 6.097033e-05, 0.0002449627, 0.0005221736, 0.001107285, 0.001107285, 
    0.0005221736, 0.0002449627, 6.097033e-05, 0,
  0, 0, 0, 0.0001398786, 0.0002967776, 0.0002967776, 0.0001398786, 0, 0, 0,
  0, 0, 0, 6.837722e-05, 0.0001459119, 0.0001459119, 6.837722e-05, 0, 0, 0,
  0, 3.013686e-05, 0.0001207906, 0.0002552228, 0.000544467, 0.000544467, 
    0.0002552228, 0.0001207906, 3.013686e-05, 0,
  0, 0.0001207906, 0.0004836885, 0.001692397, 0.001532938, 0.001532938, 
    0.001692397, 0.0004836885, 0.0001207906, 0,
  6.837722e-05, 0.0002552228, 0.001692397, 0.0009094592, 0.0003371949, 
    0.0003371949, 0.0009094592, 0.001692397, 0.0002552228, 6.837722e-05,
  0.0001459119, 0.000544467, 0.001532938, 0.0003371949, 2.186664e-05, 
    2.186664e-05, 0.0003371949, 0.001532938, 0.000544467, 0.0001459119,
  0.0001459119, 0.000544467, 0.001532938, 0.0003371949, 2.186664e-05, 
    2.186664e-05, 0.0003371949, 0.001532938, 0.000544467, 0.0001459119,
  6.837722e-05, 0.0002552228, 0.001692397, 0.0009094592, 0.0003371949, 
    0.0003371949, 0.0009094592, 0.001692397, 0.0002552228, 6.837722e-05,
  0, 0.0001207906, 0.0004836885, 0.001692397, 0.001532938, 0.001532938, 
    0.001692397, 0.0004836885, 0.0001207906, 0,
  0, 3.013686e-05, 0.0001207906, 0.0002552228, 0.000544467, 0.000544467, 
    0.0002552228, 0.0001207906, 3.013686e-05, 0,
  0, 0, 0, 6.837722e-05, 0.0001459119, 0.0001459119, 6.837722e-05, 0, 0, 0,
  0, 0, 0, 5.875934e-09, 7.011187e-09, 7.011187e-09, 5.875934e-09, 0, 0, 0,
  0, 3.286117e-09, 6.265565e-09, 2.433915e-08, 2.882667e-08, 2.882667e-08, 
    2.433915e-08, 6.265565e-09, 3.286117e-09, 0,
  0, 6.265565e-09, 2.658575e-08, 2.87517e-08, 2.54898e-08, 2.54898e-08, 
    2.87517e-08, 2.658575e-08, 6.265565e-09, 0,
  5.875934e-09, 2.433915e-08, 2.87517e-08, 2.13209e-08, 1.623442e-08, 
    1.623442e-08, 2.13209e-08, 2.87517e-08, 2.433915e-08, 5.875934e-09,
  7.011187e-09, 2.882667e-08, 2.54898e-08, 1.623442e-08, 8.385316e-09, 
    8.385316e-09, 1.623442e-08, 2.54898e-08, 2.882667e-08, 7.011187e-09,
  7.011187e-09, 2.882667e-08, 2.54898e-08, 1.623442e-08, 8.385316e-09, 
    8.385316e-09, 1.623442e-08, 2.54898e-08, 2.882667e-08, 7.011187e-09,
  5.875934e-09, 2.433915e-08, 2.87517e-08, 2.13209e-08, 1.623442e-08, 
    1.623442e-08, 2.13209e-08, 2.87517e-08, 2.433915e-08, 5.875934e-09,
  0, 6.265565e-09, 2.658575e-08, 2.87517e-08, 2.54898e-08, 2.54898e-08, 
    2.87517e-08, 2.658575e-08, 6.265565e-09, 0,
  0, 3.286117e-09, 6.265565e-09, 2.433915e-08, 2.882667e-08, 2.882667e-08, 
    2.433915e-08, 6.265565e-09, 3.286117e-09, 0,
  0, 0, 0, 5.875934e-09, 7.011187e-09, 7.011187e-09, 5.875934e-09, 0, 0, 0 ;

 vvel =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0008256877, -0.01155192, -0.0525986, -0.0525986, -0.01155192, 
    0.0008256877, 0, 0,
  0, -0.0003132102, -0.008360734, -0.00988832, -0.01105339, -0.01105339, 
    -0.00988832, -0.008360734, -0.0003132102, 0,
  0, -0.003165813, -0.005990916, -0.004564836, -0.002173914, -0.002173914, 
    -0.004564836, -0.005990916, -0.003165813, 0,
  0, -0.003779339, -0.002186223, -0.0007603604, -0.0001664206, -0.0001664206, 
    -0.0007603604, -0.002186223, -0.003779339, 0,
  0, 0.003779339, 0.002186223, 0.0007603604, 0.0001664206, 0.0001664206, 
    0.0007603604, 0.002186223, 0.003779339, 0,
  0, 0.003165813, 0.005990916, 0.004564836, 0.002173914, 0.002173914, 
    0.004564836, 0.005990916, 0.003165813, 0,
  0, 0.0003132102, 0.008360734, 0.00988832, 0.01105339, 0.01105339, 
    0.00988832, 0.008360734, 0.0003132102, 0,
  0, 0, -0.0008256877, 0.01155192, 0.0525986, 0.0525986, 0.01155192, 
    -0.0008256877, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0008988078, -0.01142125, -0.05188848, -0.05188848, -0.01142125, 
    0.0008988078, 0, 0,
  0, -0.000247678, -0.008286852, -0.009812617, -0.01079278, -0.01079278, 
    -0.009812617, -0.008286852, -0.000247678, 0,
  0, -0.003127966, -0.005943459, -0.004470771, -0.002120323, -0.002120323, 
    -0.004470771, -0.005943459, -0.003127966, 0,
  0, -0.003727764, -0.002137286, -0.000737313, -0.0001542805, -0.0001542805, 
    -0.000737313, -0.002137286, -0.003727764, 0,
  0, 0.003727764, 0.002137286, 0.000737313, 0.0001542805, 0.0001542805, 
    0.000737313, 0.002137286, 0.003727764, 0,
  0, 0.003127966, 0.005943459, 0.004470771, 0.002120323, 0.002120323, 
    0.004470771, 0.005943459, 0.003127966, 0,
  0, 0.000247678, 0.008286852, 0.009812617, 0.01079278, 0.01079278, 
    0.009812617, 0.008286852, 0.000247678, 0,
  0, 0, -0.0008988078, 0.01142125, 0.05188848, 0.05188848, 0.01142125, 
    -0.0008988078, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.001005922, -0.01098942, -0.04981515, -0.04981515, -0.01098942, 
    0.001005922, 0, 0,
  0, -0.0001338964, -0.008015784, -0.00950125, -0.01007572, -0.01007572, 
    -0.00950125, -0.008015784, -0.0001338964, 0,
  0, -0.003009181, -0.005748612, -0.004218965, -0.001982236, -0.001982236, 
    -0.004218965, -0.005748612, -0.003009181, 0,
  0, -0.00357941, -0.001999517, -0.000681401, -0.0001292175, -0.0001292175, 
    -0.000681401, -0.001999517, -0.00357941, 0,
  0, 0.00357941, 0.001999517, 0.000681401, 0.0001292175, 0.0001292175, 
    0.000681401, 0.001999517, 0.00357941, 0,
  0, 0.003009181, 0.005748612, 0.004218965, 0.001982236, 0.001982236, 
    0.004218965, 0.005748612, 0.003009181, 0,
  0, 0.0001338964, 0.008015784, 0.00950125, 0.01007572, 0.01007572, 
    0.00950125, 0.008015784, 0.0001338964, 0,
  0, 0, -0.001005922, 0.01098942, 0.04981515, 0.04981515, 0.01098942, 
    -0.001005922, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.001032454, -0.01008927, -0.04598061, -0.04598061, -0.01008927, 
    0.001032454, 0, 0,
  0, -4.092442e-05, -0.007404672, -0.00879538, -0.009030757, -0.009030757, 
    -0.00879538, -0.007404672, -4.092442e-05, 0,
  0, -0.002763917, -0.005318087, -0.003830721, -0.001783949, -0.001783949, 
    -0.003830721, -0.005318087, -0.002763917, 0,
  0, -0.003310581, -0.001799537, -0.0006064072, -0.0001023342, -0.0001023342, 
    -0.0006064072, -0.001799537, -0.003310581, 0,
  0, 0.003310581, 0.001799537, 0.0006064072, 0.0001023342, 0.0001023342, 
    0.0006064072, 0.001799537, 0.003310581, 0,
  0, 0.002763917, 0.005318087, 0.003830721, 0.001783949, 0.001783949, 
    0.003830721, 0.005318087, 0.002763917, 0,
  0, 4.092442e-05, 0.007404672, 0.00879538, 0.009030757, 0.009030757, 
    0.00879538, 0.007404672, 4.092442e-05, 0,
  0, 0, -0.001032454, 0.01008927, 0.04598061, 0.04598061, 0.01008927, 
    -0.001032454, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0009651849, -0.008752258, -0.04026955, -0.04026955, -0.008752258, 
    0.0009651849, 0, 0,
  0, 1.882779e-05, -0.006466162, -0.007693929, -0.00771859, -0.00771859, 
    -0.007693929, -0.006466162, 1.882779e-05, 0,
  0, -0.002400004, -0.004651948, -0.003310903, -0.001535694, -0.001535694, 
    -0.003310903, -0.004651948, -0.002400004, 0,
  0, -0.002906606, -0.001546011, -0.0005176318, -7.849183e-05, -7.849183e-05, 
    -0.0005176318, -0.001546011, -0.002906606, 0,
  0, 0.002906606, 0.001546011, 0.0005176318, 7.849183e-05, 7.849183e-05, 
    0.0005176318, 0.001546011, 0.002906606, 0,
  0, 0.002400004, 0.004651948, 0.003310903, 0.001535694, 0.001535694, 
    0.003310903, 0.004651948, 0.002400004, 0,
  0, -1.882779e-05, 0.006466162, 0.007693929, 0.00771859, 0.00771859, 
    0.007693929, 0.006466162, -1.882779e-05, 0,
  0, 0, -0.0009651849, 0.008752258, 0.04026955, 0.04026955, 0.008752258, 
    -0.0009651849, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0008288237, -0.007124439, -0.03311698, -0.03311698, -0.007124439, 
    0.0008288237, 0, 0,
  0, 5.001188e-05, -0.005296842, -0.006310518, -0.006221511, -0.006221511, 
    -0.006310518, -0.005296842, 5.001188e-05, 0,
  0, -0.001955896, -0.003816402, -0.002694009, -0.001249252, -0.001249252, 
    -0.002694009, -0.003816402, -0.001955896, 0,
  0, -0.002395972, -0.001252671, -0.0004183753, -5.834021e-05, -5.834021e-05, 
    -0.0004183753, -0.001252671, -0.002395972, 0,
  0, 0.002395972, 0.001252671, 0.0004183753, 5.834021e-05, 5.834021e-05, 
    0.0004183753, 0.001252671, 0.002395972, 0,
  0, 0.001955896, 0.003816402, 0.002694009, 0.001249252, 0.001249252, 
    0.002694009, 0.003816402, 0.001955896, 0,
  0, -5.001188e-05, 0.005296842, 0.006310518, 0.006221511, 0.006221511, 
    0.006310518, 0.005296842, -5.001188e-05, 0,
  0, 0, -0.0008288237, 0.007124439, 0.03311698, 0.03311698, 0.007124439, 
    -0.0008288237, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0006475092, -0.00534637, -0.02509051, -0.02509051, -0.00534637, 
    0.0006475092, 0, 0,
  0, 5.845296e-05, -0.003997323, -0.004766757, -0.004635514, -0.004635514, 
    -0.004766757, -0.003997323, 5.845296e-05, 0,
  0, -0.001469448, -0.002883687, -0.002023412, -0.000939752, -0.000939752, 
    -0.002023412, -0.002883687, -0.001469448, 0,
  0, -0.001819022, -0.0009378714, -0.0003130873, -4.102458e-05, 
    -4.102458e-05, -0.0003130873, -0.0009378714, -0.001819022, 0,
  0, 0.001819022, 0.0009378714, 0.0003130873, 4.102458e-05, 4.102458e-05, 
    0.0003130873, 0.0009378714, 0.001819022, 0,
  0, 0.001469448, 0.002883687, 0.002023412, 0.000939752, 0.000939752, 
    0.002023412, 0.002883687, 0.001469448, 0,
  0, -5.845296e-05, 0.003997323, 0.004766757, 0.004635514, 0.004635514, 
    0.004766757, 0.003997323, -5.845296e-05, 0,
  0, 0, -0.0006475092, 0.00534637, 0.02509051, 0.02509051, 0.00534637, 
    -0.0006475092, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0004403218, -0.003523594, -0.01667722, -0.01667722, -0.003523594, 
    0.0004403218, 0, 0,
  0, 4.978968e-05, -0.002647395, -0.003159238, -0.003038258, -0.003038258, 
    -0.003159238, -0.002647395, 4.978968e-05, 0,
  0, -0.0009694969, -0.001911809, -0.00133532, -0.0006215644, -0.0006215644, 
    -0.00133532, -0.001911809, -0.0009694969, 0,
  0, -0.001211213, -0.0006173779, -0.0002061807, -2.578999e-05, 
    -2.578999e-05, -0.0002061807, -0.0006173779, -0.001211213, 0,
  0, 0.001211213, 0.0006173779, 0.0002061807, 2.578999e-05, 2.578999e-05, 
    0.0002061807, 0.0006173779, 0.001211213, 0,
  0, 0.0009694969, 0.001911809, 0.00133532, 0.0006215644, 0.0006215644, 
    0.00133532, 0.001911809, 0.0009694969, 0,
  0, -4.978968e-05, 0.002647395, 0.003159238, 0.003038258, 0.003038258, 
    0.003159238, 0.002647395, -4.978968e-05, 0,
  0, 0, -0.0004403218, 0.003523594, 0.01667722, 0.01667722, 0.003523594, 
    -0.0004403218, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0002212498, -0.001726917, -0.008234199, -0.008234199, -0.001726917, 
    0.0002212498, 0, 0,
  0, 2.896606e-05, -0.001302959, -0.001555736, -0.001482464, -0.001482464, 
    -0.001555736, -0.001302959, 2.896606e-05, 0,
  0, -0.0004756116, -0.0009417262, -0.000655379, -0.0003057959, 
    -0.0003057959, -0.000655379, -0.0009417262, -0.0004756116, 0,
  0, -0.0005989244, -0.0003023877, -0.0001010627, -1.220087e-05, 
    -1.220087e-05, -0.0001010627, -0.0003023877, -0.0005989244, 0,
  0, 0.0005989244, 0.0003023877, 0.0001010627, 1.220087e-05, 1.220087e-05, 
    0.0001010627, 0.0003023877, 0.0005989244, 0,
  0, 0.0004756116, 0.0009417262, 0.000655379, 0.0003057959, 0.0003057959, 
    0.000655379, 0.0009417262, 0.0004756116, 0,
  0, -2.896606e-05, 0.001302959, 0.001555736, 0.001482464, 0.001482464, 
    0.001555736, 0.001302959, -2.896606e-05, 0,
  0, 0, -0.0002212498, 0.001726917, 0.008234199, 0.008234199, 0.001726917, 
    -0.0002212498, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -1.179029e-08, -3.384802e-08, -5.10667e-08, -5.10667e-08, 
    -3.384802e-08, -1.179029e-08, 0, 0,
  0, -1.242242e-08, -2.355311e-08, -2.524052e-08, -2.730837e-08, 
    -2.730837e-08, -2.524052e-08, -2.355311e-08, -1.242242e-08, 0,
  0, -7.061802e-09, -1.515827e-08, -1.557322e-08, -1.478742e-08, 
    -1.478742e-08, -1.557322e-08, -1.515827e-08, -7.061802e-09, 0,
  0, -2.447388e-09, -4.68496e-09, -5.164675e-09, -5.859598e-09, 
    -5.859598e-09, -5.164675e-09, -4.68496e-09, -2.447388e-09, 0,
  0, 2.447388e-09, 4.68496e-09, 5.164675e-09, 5.859598e-09, 5.859598e-09, 
    5.164675e-09, 4.68496e-09, 2.447388e-09, 0,
  0, 7.061802e-09, 1.515827e-08, 1.557322e-08, 1.478742e-08, 1.478742e-08, 
    1.557322e-08, 1.515827e-08, 7.061802e-09, 0,
  0, 1.242242e-08, 2.355311e-08, 2.524052e-08, 2.730837e-08, 2.730837e-08, 
    2.524052e-08, 2.355311e-08, 1.242242e-08, 0,
  0, 0, 1.179029e-08, 3.384802e-08, 5.10667e-08, 5.10667e-08, 3.384802e-08, 
    1.179029e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002904966, 0.002904966, 0, 0, 0, 0,
  0, 0, 0.001588732, -0.01383611, -0.01093761, -0.01093761, -0.01383611, 
    0.001588732, 0, 0,
  0, -0.0004603508, -0.008342631, -0.00982201, -0.01079595, -0.01079595, 
    -0.00982201, -0.008342631, -0.0004603508, 0,
  0, -0.002767604, -0.006091888, -0.004516106, -0.002305073, -0.002305073, 
    -0.004516106, -0.006091888, -0.002767604, 0,
  0.0001409117, -0.0005696231, -0.002037874, -0.0008045277, -0.0001358764, 
    -0.0001358764, -0.0008045277, -0.002037874, -0.0005696231, 0.0001409117,
  -0.0001409117, 0.0005696231, 0.002037874, 0.0008045277, 0.0001358764, 
    0.0001358764, 0.0008045277, 0.002037874, 0.0005696231, -0.0001409117,
  0, 0.002767604, 0.006091888, 0.004516106, 0.002305073, 0.002305073, 
    0.004516106, 0.006091888, 0.002767604, 0,
  0, 0.0004603508, 0.008342631, 0.00982201, 0.01079595, 0.01079595, 
    0.00982201, 0.008342631, 0.0004603508, 0,
  0, 0, -0.001588732, 0.01383611, 0.01093761, 0.01093761, 0.01383611, 
    -0.001588732, 0, 0,
  0, 0, 0, 0, -0.002904966, -0.002904966, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002900456, 0.002900456, 0, 0, 0, 0,
  0, 0, 0.001689613, -0.01374504, -0.01086727, -0.01086727, -0.01374504, 
    0.001689613, 0, 0,
  0, -0.0003771874, -0.008274466, -0.009729467, -0.01069149, -0.01069149, 
    -0.009729467, -0.008274466, -0.0003771874, 0,
  0, -0.002750773, -0.006040138, -0.004426829, -0.002220682, -0.002220682, 
    -0.004426829, -0.006040138, -0.002750773, 0,
  0.0001418827, -0.0005671459, -0.002014322, -0.0007758784, -0.0001304481, 
    -0.0001304481, -0.0007758784, -0.002014322, -0.0005671459, 0.0001418827,
  -0.0001418827, 0.0005671459, 0.002014322, 0.0007758784, 0.0001304481, 
    0.0001304481, 0.0007758784, 0.002014322, 0.0005671459, -0.0001418827,
  0, 0.002750773, 0.006040138, 0.004426829, 0.002220682, 0.002220682, 
    0.004426829, 0.006040138, 0.002750773, 0,
  0, 0.0003771874, 0.008274466, 0.009729467, 0.01069149, 0.01069149, 
    0.009729467, 0.008274466, 0.0003771874, 0,
  0, 0, -0.001689613, 0.01374504, 0.01086727, 0.01086727, 0.01374504, 
    -0.001689613, 0, 0,
  0, 0, 0, 0, -0.002900456, -0.002900456, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002809787, 0.002809787, 0, 0, 0, 0,
  0, 0, 0.001813428, -0.01332963, -0.01050294, -0.01050294, -0.01332963, 
    0.001813428, 0, 0,
  0, -0.0002335275, -0.008012175, -0.009390969, -0.01026892, -0.01026892, 
    -0.009390969, -0.008012175, -0.0002335275, 0,
  0, -0.00267804, -0.005836438, -0.004183661, -0.002026674, -0.002026674, 
    -0.004183661, -0.005836438, -0.00267804, 0,
  0.0001375639, -0.0005429088, -0.001930867, -0.0007077734, -0.000116664, 
    -0.000116664, -0.0007077734, -0.001930867, -0.0005429088, 0.0001375639,
  -0.0001375639, 0.0005429088, 0.001930867, 0.0007077734, 0.000116664, 
    0.000116664, 0.0007077734, 0.001930867, 0.0005429088, -0.0001375639,
  0, 0.00267804, 0.005836438, 0.004183661, 0.002026674, 0.002026674, 
    0.004183661, 0.005836438, 0.00267804, 0,
  0, 0.0002335275, 0.008012175, 0.009390969, 0.01026892, 0.01026892, 
    0.009390969, 0.008012175, 0.0002335275, 0,
  0, 0, -0.001813428, 0.01332963, 0.01050294, 0.01050294, 0.01332963, 
    -0.001813428, 0, 0,
  0, 0, 0, 0, -0.002809787, -0.002809787, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002591708, 0.002591708, 0, 0, 0, 0,
  0, 0, 0.001808339, -0.01232277, -0.009678153, -0.009678153, -0.01232277, 
    0.001808339, 0, 0,
  0, -0.0001143945, -0.007412508, -0.008663377, -0.009446746, -0.009446746, 
    -0.008663377, -0.007412508, -0.0001143945, 0,
  0, -0.002484142, -0.005389567, -0.003806251, -0.001783908, -0.001783908, 
    -0.003806251, -0.005389567, -0.002484142, 0,
  0.0001255195, -0.00049014, -0.001774436, -0.0006214951, -9.855127e-05, 
    -9.855127e-05, -0.0006214951, -0.001774436, -0.00049014, 0.0001255195,
  -0.0001255195, 0.00049014, 0.001774436, 0.0006214951, 9.855127e-05, 
    9.855127e-05, 0.0006214951, 0.001774436, 0.00049014, -0.0001255195,
  0, 0.002484142, 0.005389567, 0.003806251, 0.001783908, 0.001783908, 
    0.003806251, 0.005389567, 0.002484142, 0,
  0, 0.0001143945, 0.007412508, 0.008663377, 0.009446746, 0.009446746, 
    0.008663377, 0.007412508, 0.0001143945, 0,
  0, 0, -0.001808339, 0.01232277, 0.009678153, 0.009678153, 0.01232277, 
    -0.001808339, 0, 0,
  0, 0, 0, 0, -0.002591708, -0.002591708, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002257105, 0.002257105, 0, 0, 0, 0,
  0, 0, 0.001664641, -0.01076163, -0.008424691, -0.008424691, -0.01076163, 
    0.001664641, 0, 0,
  0, -3.382427e-05, -0.006482529, -0.007557421, -0.008239493, -0.008239493, 
    -0.007557421, -0.006482529, -3.382427e-05, 0,
  0, -0.002175087, -0.004706029, -0.003295617, -0.001509017, -0.001509017, 
    -0.003295617, -0.004706029, -0.002175087, 0,
  0.000107753, -0.0004169835, -0.001546509, -0.0005249813, -7.993602e-05, 
    -7.993602e-05, -0.0005249813, -0.001546509, -0.0004169835, 0.000107753,
  -0.000107753, 0.0004169835, 0.001546509, 0.0005249813, 7.993602e-05, 
    7.993602e-05, 0.0005249813, 0.001546509, 0.0004169835, -0.000107753,
  0, 0.002175087, 0.004706029, 0.003295617, 0.001509017, 0.001509017, 
    0.003295617, 0.004706029, 0.002175087, 0,
  0, 3.382427e-05, 0.006482529, 0.007557421, 0.008239493, 0.008239493, 
    0.007557421, 0.006482529, 3.382427e-05, 0,
  0, 0, -0.001664641, 0.01076163, 0.008424691, 0.008424691, 0.01076163, 
    -0.001664641, 0, 0,
  0, 0, 0, 0, -0.002257105, -0.002257105, 0, 0, 0, 0,
  0, 0, 0, 0, 0.001843565, 0.001843565, 0, 0, 0, 0,
  0, 0, 0.001416857, -0.008815134, -0.006879662, -0.006879662, -0.008815134, 
    0.001416857, 0, 0,
  0, 1.36996e-05, -0.005317794, -0.006185435, -0.006750421, -0.006750421, 
    -0.006185435, -0.005317794, 1.36996e-05, 0,
  0, -0.001785389, -0.003855044, -0.0026857, -0.00121061, -0.00121061, 
    -0.0026857, -0.003855044, -0.001785389, 0,
  8.679642e-05, -0.0003332556, -0.001266169, -0.0004209878, -6.231098e-05, 
    -6.231098e-05, -0.0004209878, -0.001266169, -0.0003332556, 8.679642e-05,
  -8.679642e-05, 0.0003332556, 0.001266169, 0.0004209878, 6.231098e-05, 
    6.231098e-05, 0.0004209878, 0.001266169, 0.0003332556, -8.679642e-05,
  0, 0.001785389, 0.003855044, 0.0026857, 0.00121061, 0.00121061, 0.0026857, 
    0.003855044, 0.001785389, 0,
  0, -1.36996e-05, 0.005317794, 0.006185435, 0.006750421, 0.006750421, 
    0.006185435, 0.005317794, -1.36996e-05, 0,
  0, 0, -0.001416857, 0.008815134, 0.006879662, 0.006879662, 0.008815134, 
    -0.001416857, 0, 0,
  0, 0, 0, 0, -0.001843565, -0.001843565, 0, 0, 0, 0,
  0, 0, 0, 0, 0.00138761, 0.00138761, 0, 0, 0, 0,
  0, 0, 0.001100926, -0.00665365, -0.00517776, -0.00517776, -0.00665365, 
    0.001100926, 0, 0,
  0, 3.488674e-05, -0.004019278, -0.004665238, -0.005098342, -0.005098342, 
    -0.004665238, -0.004019278, 3.488674e-05, 0,
  0, -0.001349935, -0.0029098, -0.002020023, -0.0009005336, -0.0009005336, 
    -0.002020023, -0.0029098, -0.001349935, 0,
  6.454564e-05, -0.0002460758, -0.0009557179, -0.0003131764, -4.56211e-05, 
    -4.56211e-05, -0.0003131764, -0.0009557179, -0.0002460758, 6.454564e-05,
  -6.454564e-05, 0.0002460758, 0.0009557179, 0.0003131764, 4.56211e-05, 
    4.56211e-05, 0.0003131764, 0.0009557179, 0.0002460758, -6.454564e-05,
  0, 0.001349935, 0.0029098, 0.002020023, 0.0009005336, 0.0009005336, 
    0.002020023, 0.0029098, 0.001349935, 0,
  0, -3.488674e-05, 0.004019278, 0.004665238, 0.005098342, 0.005098342, 
    0.004665238, 0.004019278, -3.488674e-05, 0,
  0, 0, -0.001100926, 0.00665365, 0.00517776, 0.00517776, 0.00665365, 
    -0.001100926, 0, 0,
  0, 0, 0, 0, -0.00138761, -0.00138761, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0009171122, 0.0009171122, 0, 0, 0, 0,
  0, 0, 0.0007463105, -0.004410344, -0.003422141, -0.003422141, -0.004410344, 
    0.0007463105, 0, 0,
  0, 3.609539e-05, -0.002667287, -0.003089655, -0.003381234, -0.003381234, 
    -0.003089655, -0.002667287, 3.609539e-05, 0,
  0, -0.0008961188, -0.001928339, -0.001335082, -0.0005902908, -0.0005902908, 
    -0.001335082, -0.001928339, -0.0008961188, 0,
  4.223891e-05, -0.0001599589, -0.0006334924, -0.0002053431, -2.968416e-05, 
    -2.968416e-05, -0.0002053431, -0.0006334924, -0.0001599589, 4.223891e-05,
  -4.223891e-05, 0.0001599589, 0.0006334924, 0.0002053431, 2.968416e-05, 
    2.968416e-05, 0.0002053431, 0.0006334924, 0.0001599589, -4.223891e-05,
  0, 0.0008961188, 0.001928339, 0.001335082, 0.0005902908, 0.0005902908, 
    0.001335082, 0.001928339, 0.0008961188, 0,
  0, -3.609539e-05, 0.002667287, 0.003089655, 0.003381234, 0.003381234, 
    0.003089655, 0.002667287, -3.609539e-05, 0,
  0, 0, -0.0007463105, 0.004410344, 0.003422141, 0.003422141, 0.004410344, 
    -0.0007463105, 0, 0,
  0, 0, 0, 0, -0.0009171122, -0.0009171122, 0, 0, 0, 0,
  0, 0, 0, 0, 0.000450985, 0.000450985, 0, 0, 0, 0,
  0, 0, 0.000374839, -0.002176257, -0.001682918, -0.001682918, -0.002176257, 
    0.000374839, 0, 0,
  0, 2.297726e-05, -0.001317347, -0.001522762, -0.001668764, -0.001668764, 
    -0.001522762, -0.001317347, 2.297726e-05, 0,
  0, -0.0004427537, -0.0009509482, -0.000656846, -0.0002885073, 
    -0.0002885073, -0.000656846, -0.0009509482, -0.0004427537, 0,
  2.061441e-05, -7.752377e-05, -0.0003124892, -0.0001004071, -1.447968e-05, 
    -1.447968e-05, -0.0001004071, -0.0003124892, -7.752377e-05, 2.061441e-05,
  -2.061441e-05, 7.752377e-05, 0.0003124892, 0.0001004071, 1.447968e-05, 
    1.447968e-05, 0.0001004071, 0.0003124892, 7.752377e-05, -2.061441e-05,
  0, 0.0004427537, 0.0009509482, 0.000656846, 0.0002885073, 0.0002885073, 
    0.000656846, 0.0009509482, 0.0004427537, 0,
  0, -2.297726e-05, 0.001317347, 0.001522762, 0.001668764, 0.001668764, 
    0.001522762, 0.001317347, -2.297726e-05, 0,
  0, 0, -0.000374839, 0.002176257, 0.001682918, 0.001682918, 0.002176257, 
    -0.000374839, 0, 0,
  0, 0, 0, 0, -0.000450985, -0.000450985, 0, 0, 0, 0,
  0, 0, 0, 0, 8.236872e-09, 8.236872e-09, 0, 0, 0, 0,
  0, 0, -1.173665e-08, -3.397699e-08, -3.650524e-08, -3.650524e-08, 
    -3.397699e-08, -1.173665e-08, 0, 0,
  0, -1.267312e-08, -2.343477e-08, -2.529044e-08, -2.602708e-08, 
    -2.602708e-08, -2.529044e-08, -2.343477e-08, -1.267312e-08, 0,
  0, -6.30858e-09, -1.545185e-08, -1.544368e-08, -1.528052e-08, 
    -1.528052e-08, -1.544368e-08, -1.545185e-08, -6.30858e-09, 0,
  -3.758351e-10, -2.031621e-09, -4.982604e-09, -5.082978e-09, -5.71314e-09, 
    -5.71314e-09, -5.082978e-09, -4.982604e-09, -2.031621e-09, -3.758351e-10,
  3.758351e-10, 2.031621e-09, 4.982604e-09, 5.082978e-09, 5.71314e-09, 
    5.71314e-09, 5.082978e-09, 4.982604e-09, 2.031621e-09, 3.758351e-10,
  0, 6.30858e-09, 1.545185e-08, 1.544368e-08, 1.528052e-08, 1.528052e-08, 
    1.544368e-08, 1.545185e-08, 6.30858e-09, 0,
  0, 1.267312e-08, 2.343477e-08, 2.529044e-08, 2.602708e-08, 2.602708e-08, 
    2.529044e-08, 2.343477e-08, 1.267312e-08, 0,
  0, 0, 1.173665e-08, 3.397699e-08, 3.650524e-08, 3.650524e-08, 3.397699e-08, 
    1.173665e-08, 0, 0,
  0, 0, 0, 0, -8.236872e-09, -8.236872e-09, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002907086, 0.002907086, 0, 0, 0, 0,
  0, 0, 0.001573083, -0.01385412, -0.01094661, -0.01094661, -0.01385412, 
    0.001573083, 0, 0,
  0, -0.0004718868, -0.008346623, -0.009787603, -0.01073877, -0.01073877, 
    -0.009787603, -0.008346623, -0.0004718868, 0,
  0, -0.002775271, -0.006071293, -0.004500326, -0.002313738, -0.002313738, 
    -0.004500326, -0.006071293, -0.002775271, 0,
  0.000141204, -0.0005710098, -0.002029181, -0.0008072912, -0.0001384091, 
    -0.0001384091, -0.0008072912, -0.002029181, -0.0005710098, 0.000141204,
  -0.000141204, 0.0005710098, 0.002029181, 0.0008072912, 0.0001384091, 
    0.0001384091, 0.0008072912, 0.002029181, 0.0005710098, -0.000141204,
  0, 0.002775271, 0.006071293, 0.004500326, 0.002313738, 0.002313738, 
    0.004500326, 0.006071293, 0.002775271, 0,
  0, 0.0004718868, 0.008346623, 0.009787603, 0.01073877, 0.01073877, 
    0.009787603, 0.008346623, 0.0004718868, 0,
  0, 0, -0.001573083, 0.01385412, 0.01094661, 0.01094661, 0.01385412, 
    -0.001573083, 0, 0,
  0, 0, 0, 0, -0.002907086, -0.002907086, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002902497, 0.002902497, 0, 0, 0, 0,
  0, 0, 0.001673691, -0.01376272, -0.01087582, -0.01087582, -0.01376272, 
    0.001673691, 0, 0,
  0, -0.000388854, -0.008278607, -0.00969515, -0.01063459, -0.01063459, 
    -0.00969515, -0.008278607, -0.000388854, 0,
  0, -0.002758372, -0.006019558, -0.004411527, -0.002229519, -0.002229519, 
    -0.004411527, -0.006019558, -0.002758372, 0,
  0.0001421608, -0.0005684611, -0.00200568, -0.0007787212, -0.0001328241, 
    -0.0001328241, -0.0007787212, -0.00200568, -0.0005684611, 0.0001421608,
  -0.0001421608, 0.0005684611, 0.00200568, 0.0007787212, 0.0001328241, 
    0.0001328241, 0.0007787212, 0.00200568, 0.0005684611, -0.0001421608,
  0, 0.002758372, 0.006019558, 0.004411527, 0.002229519, 0.002229519, 
    0.004411527, 0.006019558, 0.002758372, 0,
  0, 0.000388854, 0.008278607, 0.00969515, 0.01063459, 0.01063459, 
    0.00969515, 0.008278607, 0.000388854, 0,
  0, 0, -0.001673691, 0.01376272, 0.01087582, 0.01087582, 0.01376272, 
    -0.001673691, 0, 0,
  0, 0, 0, 0, -0.002902497, -0.002902497, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002811883, 0.002811883, 0, 0, 0, 0,
  0, 0, 0.00179794, -0.01334754, -0.01051145, -0.01051145, -0.01334754, 
    0.00179794, 0, 0,
  0, -0.0002449594, -0.008016966, -0.009357425, -0.0102144, -0.0102144, 
    -0.009357425, -0.008016966, -0.0002449594, 0,
  0, -0.002685626, -0.005816287, -0.004169604, -0.002035744, -0.002035744, 
    -0.004169604, -0.005816287, -0.002685626, 0,
  0.0001378467, -0.0005441869, -0.001922676, -0.0007107307, -0.0001187086, 
    -0.0001187086, -0.0007107307, -0.001922676, -0.0005441869, 0.0001378467,
  -0.0001378467, 0.0005441869, 0.001922676, 0.0007107307, 0.0001187086, 
    0.0001187086, 0.0007107307, 0.001922676, 0.0005441869, -0.0001378467,
  0, 0.002685626, 0.005816287, 0.004169604, 0.002035744, 0.002035744, 
    0.004169604, 0.005816287, 0.002685626, 0,
  0, 0.0002449594, 0.008016966, 0.009357425, 0.0102144, 0.0102144, 
    0.009357425, 0.008016966, 0.0002449594, 0,
  0, 0, -0.00179794, 0.01334754, 0.01051145, 0.01051145, 0.01334754, 
    -0.00179794, 0, 0,
  0, 0, 0, 0, -0.002811883, -0.002811883, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002593941, 0.002593941, 0, 0, 0, 0,
  0, 0, 0.001794341, -0.01234152, -0.009686967, -0.009686967, -0.01234152, 
    0.001794341, 0, 0,
  0, -0.0001249876, -0.007418247, -0.008632522, -0.009397025, -0.009397025, 
    -0.008632522, -0.007418247, -0.0001249876, 0,
  0, -0.002491703, -0.005371028, -0.003793863, -0.001792832, -0.001792832, 
    -0.003793863, -0.005371028, -0.002491703, 0,
  0.0001258095, -0.0004913866, -0.001767041, -0.0006244552, -0.0001002306, 
    -0.0001002306, -0.0006244552, -0.001767041, -0.0004913866, 0.0001258095,
  -0.0001258095, 0.0004913866, 0.001767041, 0.0006244552, 0.0001002306, 
    0.0001002306, 0.0006244552, 0.001767041, 0.0004913866, -0.0001258095,
  0, 0.002491703, 0.005371028, 0.003793863, 0.001792832, 0.001792832, 
    0.003793863, 0.005371028, 0.002491703, 0,
  0, 0.0001249876, 0.007418247, 0.008632522, 0.009397025, 0.009397025, 
    0.008632522, 0.007418247, 0.0001249876, 0,
  0, 0, -0.001794341, 0.01234152, 0.009686967, 0.009686967, 0.01234152, 
    -0.001794341, 0, 0,
  0, 0, 0, 0, -0.002593941, -0.002593941, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002259423, 0.002259423, 0, 0, 0, 0,
  0, 0, 0.00165294, -0.01078118, -0.008433656, -0.008433656, -0.01078118, 
    0.00165294, 0, 0,
  0, -4.305307e-05, -0.006489325, -0.007531179, -0.008196944, -0.008196944, 
    -0.007531179, -0.006489325, -4.305307e-05, 0,
  0, -0.002182445, -0.00469028, -0.003285282, -0.00151723, -0.00151723, 
    -0.003285282, -0.00469028, -0.002182445, 0,
  0.0001080338, -0.0004181444, -0.001540245, -0.000527743, -8.128507e-05, 
    -8.128507e-05, -0.000527743, -0.001540245, -0.0004181444, 0.0001080338,
  -0.0001080338, 0.0004181444, 0.001540245, 0.000527743, 8.128507e-05, 
    8.128507e-05, 0.000527743, 0.001540245, 0.0004181444, -0.0001080338,
  0, 0.002182445, 0.00469028, 0.003285282, 0.00151723, 0.00151723, 
    0.003285282, 0.00469028, 0.002182445, 0,
  0, 4.305307e-05, 0.006489325, 0.007531179, 0.008196944, 0.008196944, 
    0.007531179, 0.006489325, 4.305307e-05, 0,
  0, 0, -0.00165294, 0.01078118, 0.008433656, 0.008433656, 0.01078118, 
    -0.00165294, 0, 0,
  0, 0, 0, 0, -0.002259423, -0.002259423, 0, 0, 0, 0,
  0, 0, 0, 0, 0.00184585, 0.00184585, 0, 0, 0, 0,
  0, 0, 0.00140789, -0.008835113, -0.006888379, -0.006888379, -0.008835113, 
    0.00140789, 0, 0,
  0, 6.148277e-06, -0.005325592, -0.006165193, -0.006716882, -0.006716882, 
    -0.006165193, -0.005325592, 6.148277e-06, 0,
  0, -0.001792324, -0.003842935, -0.00267771, -0.001217658, -0.001217658, 
    -0.00267771, -0.003842935, -0.001792324, 0,
  8.704685e-05, -0.0003342622, -0.001261296, -0.0004233849, -6.336612e-05, 
    -6.336612e-05, -0.0004233849, -0.001261296, -0.0003342622, 8.704685e-05,
  -8.704685e-05, 0.0003342622, 0.001261296, 0.0004233849, 6.336612e-05, 
    6.336612e-05, 0.0004233849, 0.001261296, 0.0003342622, -8.704685e-05,
  0, 0.001792324, 0.003842935, 0.00267771, 0.001217658, 0.001217658, 
    0.00267771, 0.003842935, 0.001792324, 0,
  0, -6.148277e-06, 0.005325592, 0.006165193, 0.006716882, 0.006716882, 
    0.006165193, 0.005325592, -6.148277e-06, 0,
  0, 0, -0.00140789, 0.008835113, 0.006888379, 0.006888379, 0.008835113, 
    -0.00140789, 0, 0,
  0, 0, 0, 0, -0.00184585, -0.00184585, 0, 0, 0, 0,
  0, 0, 0, 0, 0.001389731, 0.001389731, 0, 0, 0, 0,
  0, 0, 0.001094844, -0.006673533, -0.005185776, -0.005185776, -0.006673533, 
    0.001094844, 0, 0,
  0, 2.915298e-05, -0.004027885, -0.004651777, -0.005074942, -0.005074942, 
    -0.004651777, -0.004027885, 2.915298e-05, 0,
  0, -0.001356237, -0.002901813, -0.002014543, -0.0009061344, -0.0009061344, 
    -0.002014543, -0.002901813, -0.001356237, 0,
  6.474754e-05, -0.0002468703, -0.0009523921, -0.0003151065, -4.640701e-05, 
    -4.640701e-05, -0.0003151065, -0.0009523921, -0.0002468703, 6.474754e-05,
  -6.474754e-05, 0.0002468703, 0.0009523921, 0.0003151065, 4.640701e-05, 
    4.640701e-05, 0.0003151065, 0.0009523921, 0.0002468703, -6.474754e-05,
  0, 0.001356237, 0.002901813, 0.002014543, 0.0009061344, 0.0009061344, 
    0.002014543, 0.002901813, 0.001356237, 0,
  0, -2.915298e-05, 0.004027885, 0.004651777, 0.005074942, 0.005074942, 
    0.004651777, 0.004027885, -2.915298e-05, 0,
  0, 0, -0.001094844, 0.006673533, 0.005185776, 0.005185776, 0.006673533, 
    -0.001094844, 0, 0,
  0, 0, 0, 0, -0.001389731, -0.001389731, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0009189562, 0.0009189562, 0, 0, 0, 0,
  0, 0, 0.0007430961, -0.004429145, -0.003429061, -0.003429061, -0.004429145, 
    0.0007430961, 0, 0,
  0, 3.225733e-05, -0.002676153, -0.00308317, -0.003368417, -0.003368417, 
    -0.00308317, -0.002676153, 3.225733e-05, 0,
  0, -0.0009015123, -0.001924598, -0.001332187, -0.0005942997, -0.0005942997, 
    -0.001332187, -0.001924598, -0.0009015123, 0,
  4.238164e-05, -0.0001605106, -0.0006317715, -0.0002067488, -3.021932e-05, 
    -3.021932e-05, -0.0002067488, -0.0006317715, -0.0001605106, 4.238164e-05,
  -4.238164e-05, 0.0001605106, 0.0006317715, 0.0002067488, 3.021932e-05, 
    3.021932e-05, 0.0002067488, 0.0006317715, 0.0001605106, -4.238164e-05,
  0, 0.0009015123, 0.001924598, 0.001332187, 0.0005942997, 0.0005942997, 
    0.001332187, 0.001924598, 0.0009015123, 0,
  0, -3.225733e-05, 0.002676153, 0.00308317, 0.003368417, 0.003368417, 
    0.00308317, 0.002676153, -3.225733e-05, 0,
  0, 0, -0.0007430961, 0.004429145, 0.003429061, 0.003429061, 0.004429145, 
    -0.0007430961, 0, 0,
  0, 0, 0, 0, -0.0009189562, -0.0009189562, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0004523387, 0.0004523387, 0, 0, 0, 0,
  0, 0, 0.0003742031, -0.00219062, -0.001687976, -0.001687976, -0.00219062, 
    0.0003742031, 0, 0,
  0, 2.117404e-05, -0.001324471, -0.001522253, -0.001665744, -0.001665744, 
    -0.001522253, -0.001324471, 2.117404e-05, 0,
  0, -0.0004464598, -0.0009508296, -0.0006564604, -0.0002908438, 
    -0.0002908438, -0.0006564604, -0.0009508296, -0.0004464598, 0,
  2.069441e-05, -7.782724e-05, -0.000312237, -0.0001012366, -1.477318e-05, 
    -1.477318e-05, -0.0001012366, -0.000312237, -7.782724e-05, 2.069441e-05,
  -2.069441e-05, 7.782724e-05, 0.000312237, 0.0001012366, 1.477318e-05, 
    1.477318e-05, 0.0001012366, 0.000312237, 7.782724e-05, -2.069441e-05,
  0, 0.0004464598, 0.0009508296, 0.0006564604, 0.0002908438, 0.0002908438, 
    0.0006564604, 0.0009508296, 0.0004464598, 0,
  0, -2.117404e-05, 0.001324471, 0.001522253, 0.001665744, 0.001665744, 
    0.001522253, 0.001324471, -2.117404e-05, 0,
  0, 0, -0.0003742031, 0.00219062, 0.001687976, 0.001687976, 0.00219062, 
    -0.0003742031, 0, 0,
  0, 0, 0, 0, -0.0004523387, -0.0004523387, 0, 0, 0, 0,
  0, 0, 0, 0, 8.218023e-09, 8.218023e-09, 0, 0, 0, 0,
  0, 0, -1.176477e-08, -3.397442e-08, -3.649568e-08, -3.649568e-08, 
    -3.397442e-08, -1.176477e-08, 0, 0,
  0, -1.268874e-08, -2.342423e-08, -2.524942e-08, -2.59674e-08, -2.59674e-08, 
    -2.524942e-08, -2.342423e-08, -1.268874e-08, 0,
  0, -6.309733e-09, -1.542942e-08, -1.542458e-08, -1.529537e-08, 
    -1.529537e-08, -1.542458e-08, -1.542942e-08, -6.309733e-09, 0,
  -3.793572e-10, -2.031081e-09, -4.979319e-09, -5.082796e-09, -5.735643e-09, 
    -5.735643e-09, -5.082796e-09, -4.979319e-09, -2.031081e-09, -3.793572e-10,
  3.793572e-10, 2.031081e-09, 4.979319e-09, 5.082796e-09, 5.735643e-09, 
    5.735643e-09, 5.082796e-09, 4.979319e-09, 2.031081e-09, 3.793572e-10,
  0, 6.309733e-09, 1.542942e-08, 1.542458e-08, 1.529537e-08, 1.529537e-08, 
    1.542458e-08, 1.542942e-08, 6.309733e-09, 0,
  0, 1.268874e-08, 2.342423e-08, 2.524942e-08, 2.59674e-08, 2.59674e-08, 
    2.524942e-08, 2.342423e-08, 1.268874e-08, 0,
  0, 0, 1.176477e-08, 3.397442e-08, 3.649568e-08, 3.649568e-08, 3.397442e-08, 
    1.176477e-08, 0, 0,
  0, 0, 0, 0, -8.218023e-09, -8.218023e-09, 0, 0, 0, 0,
  0, 0, 0, 0.0005927979, 0.0009220587, 0.0009220587, 0.0005927979, 0, 0, 0,
  0, 0, -0.0006781258, -0.002210401, -0.003447537, -0.003447537, 
    -0.002210401, -0.0006781258, 0, 0,
  0, -0.0002436649, -0.00828121, -0.009385014, -0.009744491, -0.009744491, 
    -0.009385014, -0.00828121, -0.0002436649, 0,
  2.937466e-05, -0.0001216534, -0.005612711, -0.004610501, -0.002375761, 
    -0.002375761, -0.004610501, -0.005612711, -0.0001216534, 2.937466e-05,
  2.721521e-05, -0.0001020982, -0.001733972, -0.0008418286, -0.000137582, 
    -0.000137582, -0.0008418286, -0.001733972, -0.0001020982, 2.721521e-05,
  -2.721521e-05, 0.0001020982, 0.001733972, 0.0008418286, 0.000137582, 
    0.000137582, 0.0008418286, 0.001733972, 0.0001020982, -2.721521e-05,
  -2.937466e-05, 0.0001216534, 0.005612711, 0.004610501, 0.002375761, 
    0.002375761, 0.004610501, 0.005612711, 0.0001216534, -2.937466e-05,
  0, 0.0002436649, 0.00828121, 0.009385014, 0.009744491, 0.009744491, 
    0.009385014, 0.00828121, 0.0002436649, 0,
  0, 0, 0.0006781258, 0.002210401, 0.003447537, 0.003447537, 0.002210401, 
    0.0006781258, 0, 0,
  0, 0, 0, -0.0005927979, -0.0009220587, -0.0009220587, -0.0005927979, 0, 0, 0,
  0, 0, 0, 0.0005801168, 0.0009105077, 0.0009105077, 0.0005801168, 0, 0, 0,
  0, 0, -0.0006111048, -0.002162982, -0.00340015, -0.00340015, -0.002162982, 
    -0.0006111048, 0, 0,
  0, -0.0001997186, -0.008210798, -0.009281811, -0.009612685, -0.009612685, 
    -0.009281811, -0.008210798, -0.0001997186, 0,
  2.753662e-05, -0.0001145652, -0.005550113, -0.00453299, -0.002300074, 
    -0.002300074, -0.00453299, -0.005550113, -0.0001145652, 2.753662e-05,
  2.698793e-05, -0.000101137, -0.001709998, -0.0008118864, -0.0001294365, 
    -0.0001294365, -0.0008118864, -0.001709998, -0.000101137, 2.698793e-05,
  -2.698793e-05, 0.000101137, 0.001709998, 0.0008118864, 0.0001294365, 
    0.0001294365, 0.0008118864, 0.001709998, 0.000101137, -2.698793e-05,
  -2.753662e-05, 0.0001145652, 0.005550113, 0.00453299, 0.002300074, 
    0.002300074, 0.00453299, 0.005550113, 0.0001145652, -2.753662e-05,
  0, 0.0001997186, 0.008210798, 0.009281811, 0.009612685, 0.009612685, 
    0.009281811, 0.008210798, 0.0001997186, 0,
  0, 0, 0.0006111048, 0.002162982, 0.00340015, 0.00340015, 0.002162982, 
    0.0006111048, 0, 0,
  0, 0, 0, -0.0005801168, -0.0009105077, -0.0009105077, -0.0005801168, 0, 0, 0,
  0, 0, 0, 0.0005478773, 0.0008747906, 0.0008747906, 0.0005478773, 0, 0, 0,
  0, 0, -0.0004923516, -0.002043155, -0.003264622, -0.003264622, 
    -0.002043155, -0.0004923516, 0, 0,
  0, -0.0001212417, -0.007942389, -0.008962078, -0.009233337, -0.009233337, 
    -0.008962078, -0.007942389, -0.0001212417, 0,
  2.459871e-05, -0.0001018609, -0.005351122, -0.004296739, -0.00210894, 
    -0.00210894, -0.004296739, -0.005351122, -0.0001018609, 2.459871e-05,
  2.619718e-05, -9.80252e-05, -0.001640004, -0.0007429817, -0.0001134368, 
    -0.0001134368, -0.0007429817, -0.001640004, -9.80252e-05, 2.619718e-05,
  -2.619718e-05, 9.80252e-05, 0.001640004, 0.0007429817, 0.0001134368, 
    0.0001134368, 0.0007429817, 0.001640004, 9.80252e-05, -2.619718e-05,
  -2.459871e-05, 0.0001018609, 0.005351122, 0.004296739, 0.00210894, 
    0.00210894, 0.004296739, 0.005351122, 0.0001018609, -2.459871e-05,
  0, 0.0001212417, 0.007942389, 0.008962078, 0.009233337, 0.009233337, 
    0.008962078, 0.007942389, 0.0001212417, 0,
  0, 0, 0.0004923516, 0.002043155, 0.003264622, 0.003264622, 0.002043155, 
    0.0004923516, 0, 0,
  0, 0, 0, -0.0005478773, -0.0008747906, -0.0008747906, -0.0005478773, 0, 0, 0,
  0, 0, 0, 0.0004952688, 0.0008008862, 0.0008008862, 0.0004952688, 0, 0, 0,
  0, 0, -0.0003777269, -0.001847067, -0.002988057, -0.002988057, 
    -0.001847067, -0.0003777269, 0, 0,
  0, -5.588763e-05, -0.007337223, -0.008294187, -0.008522817, -0.008522817, 
    -0.008294187, -0.007337223, -5.588763e-05, 0,
  2.114013e-05, -8.658683e-05, -0.004942738, -0.003911743, -0.001860625, 
    -0.001860625, -0.003911743, -0.004942738, -8.658683e-05, 2.114013e-05,
  2.395063e-05, -8.959212e-05, -0.001511542, -0.0006553119, -9.445607e-05, 
    -9.445607e-05, -0.0006553119, -0.001511542, -8.959212e-05, 2.395063e-05,
  -2.395063e-05, 8.959212e-05, 0.001511542, 0.0006553119, 9.445607e-05, 
    9.445607e-05, 0.0006553119, 0.001511542, 8.959212e-05, -2.395063e-05,
  -2.114013e-05, 8.658683e-05, 0.004942738, 0.003911743, 0.001860625, 
    0.001860625, 0.003911743, 0.004942738, 8.658683e-05, -2.114013e-05,
  0, 5.588763e-05, 0.007337223, 0.008294187, 0.008522817, 0.008522817, 
    0.008294187, 0.007337223, 5.588763e-05, 0,
  0, 0, 0.0003777269, 0.001847067, 0.002988057, 0.002988057, 0.001847067, 
    0.0003777269, 0, 0,
  0, 0, 0, -0.0004952688, -0.0008008862, -0.0008008862, -0.0004952688, 0, 0, 0,
  0, 0, 0, 0.0004246696, 0.0006926283, 0.0006926283, 0.0004246696, 0, 0, 0,
  0, 0, -0.0002782268, -0.001583891, -0.002583976, -0.002583976, 
    -0.001583891, -0.0002782268, 0, 0,
  0, -1.112143e-05, -0.006408261, -0.007265355, -0.007463949, -0.007463949, 
    -0.007265355, -0.006408261, -1.112143e-05, 0,
  1.734022e-05, -7.011503e-05, -0.004321288, -0.003385333, -0.001574976, 
    -0.001574976, -0.003385333, -0.004321288, -7.011503e-05, 1.734022e-05,
  2.057202e-05, -7.694183e-05, -0.001321844, -0.0005555307, -7.596873e-05, 
    -7.596873e-05, -0.0005555307, -0.001321844, -7.694183e-05, 2.057202e-05,
  -2.057202e-05, 7.694183e-05, 0.001321844, 0.0005555307, 7.596873e-05, 
    7.596873e-05, 0.0005555307, 0.001321844, 7.694183e-05, -2.057202e-05,
  -1.734022e-05, 7.011503e-05, 0.004321288, 0.003385333, 0.001574976, 
    0.001574976, 0.003385333, 0.004321288, 7.011503e-05, -1.734022e-05,
  0, 1.112143e-05, 0.006408261, 0.007265355, 0.007463949, 0.007463949, 
    0.007265355, 0.006408261, 1.112143e-05, 0,
  0, 0, 0.0002782268, 0.001583891, 0.002583976, 0.002583976, 0.001583891, 
    0.0002782268, 0, 0,
  0, 0, 0, -0.0004246696, -0.0006926283, -0.0006926283, -0.0004246696, 0, 0, 0,
  0, 0, 0, 0.0003426427, 0.0005622989, 0.0005622989, 0.0003426427, 0, 0, 0,
  0, 0, -0.0001949756, -0.001278079, -0.002097788, -0.002097788, 
    -0.001278079, -0.0001949756, 0, 0,
  0, 1.515912e-05, -0.005252321, -0.00597164, -0.006139196, -0.006139196, 
    -0.00597164, -0.005252321, 1.515912e-05, 0,
  1.346958e-05, -5.373624e-05, -0.003545666, -0.00275675, -0.001263427, 
    -0.001263427, -0.00275675, -0.003545666, -5.373624e-05, 1.346958e-05,
  1.65724e-05, -6.196715e-05, -0.001085737, -0.0004466841, -5.899592e-05, 
    -5.899592e-05, -0.0004466841, -0.001085737, -6.196715e-05, 1.65724e-05,
  -1.65724e-05, 6.196715e-05, 0.001085737, 0.0004466841, 5.899592e-05, 
    5.899592e-05, 0.0004466841, 0.001085737, 6.196715e-05, -1.65724e-05,
  -1.346958e-05, 5.373624e-05, 0.003545666, 0.00275675, 0.001263427, 
    0.001263427, 0.00275675, 0.003545666, 5.373624e-05, -1.346958e-05,
  0, -1.515912e-05, 0.005252321, 0.00597164, 0.006139196, 0.006139196, 
    0.00597164, 0.005252321, -1.515912e-05, 0,
  0, 0, 0.0001949756, 0.001278079, 0.002097788, 0.002097788, 0.001278079, 
    0.0001949756, 0, 0,
  0, 0, 0, -0.0003426427, -0.0005622989, -0.0005622989, -0.0003426427, 0, 0, 0,
  0, 0, 0, 0.0002554594, 0.0004210924, 0.0004210924, 0.0002554594, 0, 0, 0,
  0, 0, -0.0001277715, -0.0009529833, -0.001571069, -0.001571069, 
    -0.0009529833, -0.0001277715, 0, 0,
  0, 2.597713e-05, -0.003969084, -0.004523174, -0.004654329, -0.004654329, 
    -0.004523174, -0.003969084, 2.597713e-05, 0,
  9.73296e-06, -3.829425e-05, -0.002681595, -0.002072225, -0.000939663, 
    -0.000939663, -0.002072225, -0.002681595, -3.829425e-05, 9.73296e-06,
  1.231937e-05, -4.604799e-05, -0.0008220871, -0.0003330655, -4.315929e-05, 
    -4.315929e-05, -0.0003330655, -0.0008220871, -4.604799e-05, 1.231937e-05,
  -1.231937e-05, 4.604799e-05, 0.0008220871, 0.0003330655, 4.315929e-05, 
    4.315929e-05, 0.0003330655, 0.0008220871, 4.604799e-05, -1.231937e-05,
  -9.73296e-06, 3.829425e-05, 0.002681595, 0.002072225, 0.000939663, 
    0.000939663, 0.002072225, 0.002681595, 3.829425e-05, -9.73296e-06,
  0, -2.597713e-05, 0.003969084, 0.004523174, 0.004654329, 0.004654329, 
    0.004523174, 0.003969084, -2.597713e-05, 0,
  0, 0, 0.0001277715, 0.0009529833, 0.001571069, 0.001571069, 0.0009529833, 
    0.0001277715, 0, 0,
  0, 0, 0, -0.0002554594, -0.0004210924, -0.0004210924, -0.0002554594, 0, 0, 0,
  0, 0, 0, 0.0001676652, 0.0002771921, 0.0002771921, 0.0001676652, 0, 0, 0,
  0, 0, -7.482824e-05, -0.000625542, -0.001034266, -0.001034266, 
    -0.000625542, -7.482824e-05, 0, 0,
  0, 2.485497e-05, -0.002636307, -0.003009646, -0.003099435, -0.003099435, 
    -0.003009646, -0.002636307, 2.485497e-05, 0,
  6.229418e-06, -2.415505e-05, -0.001781949, -0.001369582, -0.0006161059, 
    -0.0006161059, -0.001369582, -0.001781949, -2.415505e-05, 6.229418e-06,
  8.053987e-06, -3.009092e-05, -0.0005467999, -0.0002189408, -2.812003e-05, 
    -2.812003e-05, -0.0002189408, -0.0005467999, -3.009092e-05, 8.053987e-06,
  -8.053987e-06, 3.009092e-05, 0.0005467999, 0.0002189408, 2.812003e-05, 
    2.812003e-05, 0.0002189408, 0.0005467999, 3.009092e-05, -8.053987e-06,
  -6.229418e-06, 2.415505e-05, 0.001781949, 0.001369582, 0.0006161059, 
    0.0006161059, 0.001369582, 0.001781949, 2.415505e-05, -6.229418e-06,
  0, -2.485497e-05, 0.002636307, 0.003009646, 0.003099435, 0.003099435, 
    0.003009646, 0.002636307, -2.485497e-05, 0,
  0, 0, 7.482824e-05, 0.000625542, 0.001034266, 0.001034266, 0.000625542, 
    7.482824e-05, 0, 0,
  0, 0, 0, -0.0001676652, -0.0002771921, -0.0002771921, -0.0001676652, 0, 0, 0,
  0, 0, 0, 8.20508e-05, 0.0001358988, 0.0001358988, 8.20508e-05, 0, 0, 0,
  0, 0, -3.311473e-05, -0.0003061637, -0.0005071203, -0.0005071203, 
    -0.0003061637, -3.311473e-05, 0, 0,
  0, 1.538461e-05, -0.00130512, -0.00149255, -0.00153842, -0.00153842, 
    -0.00149255, -0.00130512, 1.538461e-05, 0,
  2.978258e-06, -1.13621e-05, -0.000882685, -0.0006751646, -0.0003017059, 
    -0.0003017059, -0.0006751646, -0.000882685, -1.13621e-05, 2.978258e-06,
  3.9232e-06, -1.464857e-05, -0.0002710968, -0.000107478, -1.377299e-05, 
    -1.377299e-05, -0.000107478, -0.0002710968, -1.464857e-05, 3.9232e-06,
  -3.9232e-06, 1.464857e-05, 0.0002710968, 0.000107478, 1.377299e-05, 
    1.377299e-05, 0.000107478, 0.0002710968, 1.464857e-05, -3.9232e-06,
  -2.978258e-06, 1.13621e-05, 0.000882685, 0.0006751646, 0.0003017059, 
    0.0003017059, 0.0006751646, 0.000882685, 1.13621e-05, -2.978258e-06,
  0, -1.538461e-05, 0.00130512, 0.00149255, 0.00153842, 0.00153842, 
    0.00149255, 0.00130512, -1.538461e-05, 0,
  0, 0, 3.311473e-05, 0.0003061637, 0.0005071203, 0.0005071203, 0.0003061637, 
    3.311473e-05, 0, 0,
  0, 0, 0, -8.20508e-05, -0.0001358988, -0.0001358988, -8.20508e-05, 0, 0, 0,
  0, 0, 0, 5.808732e-09, 7.001435e-09, 7.001435e-09, 5.808732e-09, 0, 0, 0,
  0, 0, -1.320141e-08, -2.375368e-08, -2.863566e-08, -2.863566e-08, 
    -2.375368e-08, -1.320141e-08, 0, 0,
  0, -1.151457e-08, -2.347333e-08, -2.46941e-08, -2.551781e-08, 
    -2.551781e-08, -2.46941e-08, -2.347333e-08, -1.151457e-08, 0,
  5.853413e-10, -4.234781e-09, -1.558718e-08, -1.544228e-08, -1.530671e-08, 
    -1.530671e-08, -1.544228e-08, -1.558718e-08, -4.234781e-09, 5.853413e-10,
  3.118638e-10, -1.096469e-09, -4.875147e-09, -5.093391e-09, -5.799936e-09, 
    -5.799936e-09, -5.093391e-09, -4.875147e-09, -1.096469e-09, 3.118638e-10,
  -3.118638e-10, 1.096469e-09, 4.875147e-09, 5.093391e-09, 5.799936e-09, 
    5.799936e-09, 5.093391e-09, 4.875147e-09, 1.096469e-09, -3.118638e-10,
  -5.853413e-10, 4.234781e-09, 1.558718e-08, 1.544228e-08, 1.530671e-08, 
    1.530671e-08, 1.544228e-08, 1.558718e-08, 4.234781e-09, -5.853413e-10,
  0, 1.151457e-08, 2.347333e-08, 2.46941e-08, 2.551781e-08, 2.551781e-08, 
    2.46941e-08, 2.347333e-08, 1.151457e-08, 0,
  0, 0, 1.320141e-08, 2.375368e-08, 2.863566e-08, 2.863566e-08, 2.375368e-08, 
    1.320141e-08, 0, 0,
  0, 0, 0, -5.808732e-09, -7.001435e-09, -7.001435e-09, -5.808732e-09, 0, 0, 0,
  0, 0, 0, 0.0005976551, 0.0009266008, 0.0009266008, 0.0005976551, 0, 0, 0,
  0, 0, -0.0006940318, -0.002228644, -0.00346467, -0.00346467, -0.002228644, 
    -0.0006940318, 0, 0,
  0, -0.0002546235, -0.00828829, -0.009351598, -0.009684209, -0.009684209, 
    -0.009351598, -0.00828829, -0.0002546235, 0,
  3.046667e-05, -0.0001257831, -0.005597732, -0.004594702, -0.002380941, 
    -0.002380941, -0.004594702, -0.005597732, -0.0001257831, 3.046667e-05,
  2.745757e-05, -0.00010299, -0.001725802, -0.0008440774, -0.0001401419, 
    -0.0001401419, -0.0008440774, -0.001725802, -0.00010299, 2.745757e-05,
  -2.745757e-05, 0.00010299, 0.001725802, 0.0008440774, 0.0001401419, 
    0.0001401419, 0.0008440774, 0.001725802, 0.00010299, -2.745757e-05,
  -3.046667e-05, 0.0001257831, 0.005597732, 0.004594702, 0.002380941, 
    0.002380941, 0.004594702, 0.005597732, 0.0001257831, -3.046667e-05,
  0, 0.0002546235, 0.00828829, 0.009351598, 0.009684209, 0.009684209, 
    0.009351598, 0.00828829, 0.0002546235, 0,
  0, 0, 0.0006940318, 0.002228644, 0.00346467, 0.00346467, 0.002228644, 
    0.0006940318, 0, 0,
  0, 0, 0, -0.0005976551, -0.0009266008, -0.0009266008, -0.0005976551, 0, 0, 0,
  0, 0, 0, 0.000584978, 0.0009150683, 0.0009150683, 0.000584978, 0, 0, 0,
  0, 0, -0.0006271242, -0.002181178, -0.003417269, -0.003417269, 
    -0.002181178, -0.0006271242, 0, 0,
  0, -0.0002107615, -0.008217847, -0.00924895, -0.009553849, -0.009553849, 
    -0.00924895, -0.008217847, -0.0002107615, 0,
  2.863302e-05, -0.0001186984, -0.005535415, -0.004517405, -0.002305315, 
    -0.002305315, -0.004517405, -0.005535415, -0.0001186984, 2.863302e-05,
  2.72283e-05, -0.0001020216, -0.001702062, -0.0008142332, -0.0001318761, 
    -0.0001318761, -0.0008142332, -0.001702062, -0.0001020216, 2.72283e-05,
  -2.72283e-05, 0.0001020216, 0.001702062, 0.0008142332, 0.0001318761, 
    0.0001318761, 0.0008142332, 0.001702062, 0.0001020216, -2.72283e-05,
  -2.863302e-05, 0.0001186984, 0.005535415, 0.004517405, 0.002305315, 
    0.002305315, 0.004517405, 0.005535415, 0.0001186984, -2.863302e-05,
  0, 0.0002107615, 0.008217847, 0.00924895, 0.009553849, 0.009553849, 
    0.00924895, 0.008217847, 0.0002107615, 0,
  0, 0, 0.0006271242, 0.002181178, 0.003417269, 0.003417269, 0.002181178, 
    0.0006271242, 0, 0,
  0, 0, 0, -0.000584978, -0.0009150683, -0.0009150683, -0.000584978, 0, 0, 0,
  0, 0, 0, 0.0005526862, 0.0008792863, 0.0008792863, 0.0005526862, 0, 0, 0,
  0, 0, -0.0005080745, -0.002061121, -0.00328145, -0.00328145, -0.002061121, 
    -0.0005080745, 0, 0,
  0, -0.0001321262, -0.007949643, -0.008930719, -0.009177702, -0.009177702, 
    -0.008930719, -0.007949643, -0.0001321262, 0,
  2.568198e-05, -0.0001059302, -0.005337188, -0.004282035, -0.002114474, 
    -0.002114474, -0.004282035, -0.005337188, -0.0001059302, 2.568198e-05,
  2.642871e-05, -9.887929e-05, -0.001632569, -0.000745484, -0.000115579, 
    -0.000115579, -0.000745484, -0.001632569, -9.887929e-05, 2.642871e-05,
  -2.642871e-05, 9.887929e-05, 0.001632569, 0.000745484, 0.000115579, 
    0.000115579, 0.000745484, 0.001632569, 9.887929e-05, -2.642871e-05,
  -2.568198e-05, 0.0001059302, 0.005337188, 0.004282035, 0.002114474, 
    0.002114474, 0.004282035, 0.005337188, 0.0001059302, -2.568198e-05,
  0, 0.0001321262, 0.007949643, 0.008930719, 0.009177702, 0.009177702, 
    0.008930719, 0.007949643, 0.0001321262, 0,
  0, 0, 0.0005080745, 0.002061121, 0.00328145, 0.00328145, 0.002061121, 
    0.0005080745, 0, 0,
  0, 0, 0, -0.0005526862, -0.0008792863, -0.0008792863, -0.0005526862, 0, 0, 0,
  0, 0, 0, 0.0004998034, 0.0008051077, 0.0008051077, 0.0004998034, 0, 0, 0,
  0, 0, -0.0003924186, -0.001863993, -0.003003838, -0.003003838, 
    -0.001863993, -0.0003924186, 0, 0,
  0, -6.606273e-05, -0.007344917, -0.008265833, -0.0084723, -0.0084723, 
    -0.008265833, -0.007344917, -6.606273e-05, 0,
  2.215118e-05, -9.037773e-05, -0.004930267, -0.00389852, -0.00186627, 
    -0.00186627, -0.00389852, -0.004930267, -9.037773e-05, 2.215118e-05,
  2.416347e-05, -9.037944e-05, -0.001504841, -0.0006578621, -9.625436e-05, 
    -9.625436e-05, -0.0006578621, -0.001504841, -9.037944e-05, 2.416347e-05,
  -2.416347e-05, 9.037944e-05, 0.001504841, 0.0006578621, 9.625436e-05, 
    9.625436e-05, 0.0006578621, 0.001504841, 9.037944e-05, -2.416347e-05,
  -2.215118e-05, 9.037773e-05, 0.004930267, 0.00389852, 0.00186627, 
    0.00186627, 0.00389852, 0.004930267, 9.037773e-05, -2.215118e-05,
  0, 6.606273e-05, 0.007344917, 0.008265833, 0.0084723, 0.0084723, 
    0.008265833, 0.007344917, 6.606273e-05, 0,
  0, 0, 0.0003924186, 0.001863993, 0.003003838, 0.003003838, 0.001863993, 
    0.0003924186, 0, 0,
  0, 0, 0, -0.0004998034, -0.0008051077, -0.0008051077, -0.0004998034, 0, 0, 0,
  0, 0, 0, 0.0004287128, 0.0006963831, 0.0006963831, 0.0004287128, 0, 0, 0,
  0, 0, -0.0002912104, -0.001598977, -0.002598002, -0.002598002, 
    -0.001598977, -0.0002912104, 0, 0,
  0, -2.007348e-05, -0.006416466, -0.007241611, -0.007420705, -0.007420705, 
    -0.007241611, -0.006416466, -2.007348e-05, 0,
  1.822705e-05, -7.34364e-05, -0.00431102, -0.00337412, -0.001580322, 
    -0.001580322, -0.00337412, -0.00431102, -7.34364e-05, 1.822705e-05,
  2.07577e-05, -7.763013e-05, -0.001316148, -0.0005579437, -7.744075e-05, 
    -7.744075e-05, -0.0005579437, -0.001316148, -7.763013e-05, 2.07577e-05,
  -2.07577e-05, 7.763013e-05, 0.001316148, 0.0005579437, 7.744075e-05, 
    7.744075e-05, 0.0005579437, 0.001316148, 7.763013e-05, -2.07577e-05,
  -1.822705e-05, 7.34364e-05, 0.00431102, 0.00337412, 0.001580322, 
    0.001580322, 0.00337412, 0.00431102, 7.34364e-05, -1.822705e-05,
  0, 2.007348e-05, 0.006416466, 0.007241611, 0.007420705, 0.007420705, 
    0.007241611, 0.006416466, 2.007348e-05, 0,
  0, 0, 0.0002912104, 0.001598977, 0.002598002, 0.002598002, 0.001598977, 
    0.0002912104, 0, 0,
  0, 0, 0, -0.0004287128, -0.0006963831, -0.0006963831, -0.0004287128, 0, 0, 0,
  0, 0, 0, 0.0003460448, 0.0005654459, 0.0005654459, 0.0003460448, 0, 0, 0,
  0, 0, -0.0002058307, -0.001290771, -0.002109539, -0.002109539, 
    -0.001290771, -0.0002058307, 0, 0,
  0, 7.749403e-06, -0.005260962, -0.005953672, -0.006104944, -0.006104944, 
    -0.005953672, -0.005260962, 7.749403e-06, 0,
  1.419874e-05, -5.646477e-05, -0.003538133, -0.002747942, -0.001268135, 
    -0.001268135, -0.002747942, -0.003538133, -5.646477e-05, 1.419874e-05,
  1.672446e-05, -6.253186e-05, -0.001081273, -0.000448809, -6.016145e-05, 
    -6.016145e-05, -0.000448809, -0.001081273, -6.253186e-05, 1.672446e-05,
  -1.672446e-05, 6.253186e-05, 0.001081273, 0.000448809, 6.016145e-05, 
    6.016145e-05, 0.000448809, 0.001081273, 6.253186e-05, -1.672446e-05,
  -1.419874e-05, 5.646477e-05, 0.003538133, 0.002747942, 0.001268135, 
    0.001268135, 0.002747942, 0.003538133, 5.646477e-05, -1.419874e-05,
  0, -7.749403e-06, 0.005260962, 0.005953672, 0.006104944, 0.006104944, 
    0.005953672, 0.005260962, -7.749403e-06, 0,
  0, 0, 0.0002058307, 0.001290771, 0.002109539, 0.002109539, 0.001290771, 
    0.0002058307, 0, 0,
  0, 0, 0, -0.0003460448, -0.0005654459, -0.0005654459, -0.0003460448, 0, 0, 0,
  0, 0, 0, 0.0002581271, 0.0004235449, 0.0004235449, 0.0002581271, 0, 0, 0,
  0, 0, -0.0001362561, -0.0009629345, -0.001580223, -0.001580223, 
    -0.0009629345, -0.0001362561, 0, 0,
  0, 2.028637e-05, -0.003977902, -0.004511587, -0.004630116, -0.004630116, 
    -0.004511587, -0.003977902, 2.028637e-05, 0,
  1.02857e-05, -4.036111e-05, -0.002677063, -0.002066068, -0.000943519, 
    -0.000943519, -0.002066068, -0.002677063, -4.036111e-05, 1.02857e-05,
  1.243415e-05, -4.647492e-05, -0.0008189927, -0.0003348062, -4.403178e-05, 
    -4.403178e-05, -0.0003348062, -0.0008189927, -4.647492e-05, 1.243415e-05,
  -1.243415e-05, 4.647492e-05, 0.0008189927, 0.0003348062, 4.403178e-05, 
    4.403178e-05, 0.0003348062, 0.0008189927, 4.647492e-05, -1.243415e-05,
  -1.02857e-05, 4.036111e-05, 0.002677063, 0.002066068, 0.000943519, 
    0.000943519, 0.002066068, 0.002677063, 4.036111e-05, -1.02857e-05,
  0, -2.028637e-05, 0.003977902, 0.004511587, 0.004630116, 0.004630116, 
    0.004511587, 0.003977902, -2.028637e-05, 0,
  0, 0, 0.0001362561, 0.0009629345, 0.001580223, 0.001580223, 0.0009629345, 
    0.0001362561, 0, 0,
  0, 0, 0, -0.0002581271, -0.0004235449, -0.0004235449, -0.0002581271, 0, 0, 0,
  0, 0, 0, 0.0001695268, 0.0002789027, 0.0002789027, 0.0001695268, 0, 0, 0,
  0, 0, -8.068501e-05, -0.0006324865, -0.00104065, -0.00104065, 
    -0.0006324865, -8.068501e-05, 0, 0,
  0, 2.103172e-05, -0.002644493, -0.003004336, -0.003085589, -0.003085589, 
    -0.003004336, -0.002644493, 2.103172e-05, 0,
  6.594866e-06, -2.552069e-05, -0.001780329, -0.001366226, -0.0006189904, 
    -0.0006189904, -0.001366226, -0.001780329, -2.552069e-05, 6.594866e-06,
  8.130642e-06, -3.037642e-05, -0.0005451211, -0.0002202333, -2.871067e-05, 
    -2.871067e-05, -0.0002202333, -0.0005451211, -3.037642e-05, 8.130642e-06,
  -8.130642e-06, 3.037642e-05, 0.0005451211, 0.0002202333, 2.871067e-05, 
    2.871067e-05, 0.0002202333, 0.0005451211, 3.037642e-05, -8.130642e-06,
  -6.594866e-06, 2.552069e-05, 0.001780329, 0.001366226, 0.0006189904, 
    0.0006189904, 0.001366226, 0.001780329, 2.552069e-05, -6.594866e-06,
  0, -2.103172e-05, 0.002644493, 0.003004336, 0.003085589, 0.003085589, 
    0.003004336, 0.002644493, -2.103172e-05, 0,
  0, 0, 8.068501e-05, 0.0006324865, 0.00104065, 0.00104065, 0.0006324865, 
    8.068501e-05, 0, 0,
  0, 0, 0, -0.0001695268, -0.0002789027, -0.0002789027, -0.0001695268, 0, 0, 0,
  0, 0, 0, 8.301486e-05, 0.0001368101, 0.0001368101, 8.301486e-05, 0, 0, 0,
  0, 0, -3.599225e-05, -0.0003097604, -0.0005105206, -0.0005105206, 
    -0.0003097604, -3.599225e-05, 0, 0,
  0, 1.357571e-05, -0.001310641, -0.001491929, -0.001533798, -0.001533798, 
    -0.001491929, -0.001310641, 1.357571e-05, 0,
  3.150988e-06, -1.200721e-05, -0.0008830633, -0.0006744439, -0.0003034991, 
    -0.0003034991, -0.0006744439, -0.0008830633, -1.200721e-05, 3.150988e-06,
  3.961909e-06, -1.479293e-05, -0.0002706518, -0.0001082485, -1.408372e-05, 
    -1.408372e-05, -0.0001082485, -0.0002706518, -1.479293e-05, 3.961909e-06,
  -3.961909e-06, 1.479293e-05, 0.0002706518, 0.0001082485, 1.408372e-05, 
    1.408372e-05, 0.0001082485, 0.0002706518, 1.479293e-05, -3.961909e-06,
  -3.150988e-06, 1.200721e-05, 0.0008830633, 0.0006744439, 0.0003034991, 
    0.0003034991, 0.0006744439, 0.0008830633, 1.200721e-05, -3.150988e-06,
  0, -1.357571e-05, 0.001310641, 0.001491929, 0.001533798, 0.001533798, 
    0.001491929, 0.001310641, -1.357571e-05, 0,
  0, 0, 3.599225e-05, 0.0003097604, 0.0005105206, 0.0005105206, 0.0003097604, 
    3.599225e-05, 0, 0,
  0, 0, 0, -8.301486e-05, -0.0001368101, -0.0001368101, -8.301486e-05, 0, 0, 0,
  0, 0, 0, 5.811907e-09, 7.001984e-09, 7.001984e-09, 5.811907e-09, 0, 0, 0,
  0, 0, -1.323016e-08, -2.378301e-08, -2.865949e-08, -2.865949e-08, 
    -2.378301e-08, -1.323016e-08, 0, 0,
  0, -1.152815e-08, -2.346661e-08, -2.464363e-08, -2.544626e-08, 
    -2.544626e-08, -2.464363e-08, -2.346661e-08, -1.152815e-08, 0,
  5.855569e-10, -4.240657e-09, -1.557423e-08, -1.542444e-08, -1.531423e-08, 
    -1.531423e-08, -1.542444e-08, -1.557423e-08, -4.240657e-09, 5.855569e-10,
  3.119792e-10, -1.097102e-09, -4.872368e-09, -5.09584e-09, -5.821105e-09, 
    -5.821105e-09, -5.09584e-09, -4.872368e-09, -1.097102e-09, 3.119792e-10,
  -3.119792e-10, 1.097102e-09, 4.872368e-09, 5.09584e-09, 5.821105e-09, 
    5.821105e-09, 5.09584e-09, 4.872368e-09, 1.097102e-09, -3.119792e-10,
  -5.855569e-10, 4.240657e-09, 1.557423e-08, 1.542444e-08, 1.531423e-08, 
    1.531423e-08, 1.542444e-08, 1.557423e-08, 4.240657e-09, -5.855569e-10,
  0, 1.152815e-08, 2.346661e-08, 2.464363e-08, 2.544626e-08, 2.544626e-08, 
    2.464363e-08, 2.346661e-08, 1.152815e-08, 0,
  0, 0, 1.323016e-08, 2.378301e-08, 2.865949e-08, 2.865949e-08, 2.378301e-08, 
    1.323016e-08, 0, 0,
  0, 0, 0, -5.811907e-09, -7.001984e-09, -7.001984e-09, -5.811907e-09, 0, 0, 0,
  0, 0, 0, 0.0006019049, 0.0009306039, 0.0009306039, 0.0006019049, 0, 0, 0,
  0, 0, -0.0007108127, -0.002244591, -0.003479775, -0.003479775, 
    -0.002244591, -0.0007108127, 0, 0,
  0, -0.0002657369, -0.008294973, -0.009318897, -0.009625057, -0.009625057, 
    -0.009318897, -0.008294973, -0.0002657369, 0,
  3.147144e-05, -0.0001295755, -0.005582972, -0.004578956, -0.002385959, 
    -0.002385959, -0.004578956, -0.005582972, -0.0001295755, 3.147144e-05,
  2.767998e-05, -0.0001038073, -0.001717737, -0.0008463032, -0.0001427074, 
    -0.0001427074, -0.0008463032, -0.001717737, -0.0001038073, 2.767998e-05,
  -2.767998e-05, 0.0001038073, 0.001717737, 0.0008463032, 0.0001427074, 
    0.0001427074, 0.0008463032, 0.001717737, 0.0001038073, -2.767998e-05,
  -3.147144e-05, 0.0001295755, 0.005582972, 0.004578956, 0.002385959, 
    0.002385959, 0.004578956, 0.005582972, 0.0001295755, -3.147144e-05,
  0, 0.0002657369, 0.008294973, 0.009318897, 0.009625057, 0.009625057, 
    0.009318897, 0.008294973, 0.0002657369, 0,
  0, 0, 0.0007108127, 0.002244591, 0.003479775, 0.003479775, 0.002244591, 
    0.0007108127, 0, 0,
  0, 0, 0, -0.0006019049, -0.0009306039, -0.0009306039, -0.0006019049, 0, 0, 0,
  0, 0, 0, 0.0005892332, 0.0009190909, 0.0009190909, 0.0005892332, 0, 0, 0,
  0, 0, -0.0006440201, -0.002197089, -0.00343237, -0.00343237, -0.002197089, 
    -0.0006440201, 0, 0,
  0, -0.0002219629, -0.008224508, -0.009216779, -0.009496097, -0.009496097, 
    -0.009216779, -0.008224508, -0.0002219629, 0,
  2.964231e-05, -0.0001224955, -0.005520921, -0.004501875, -0.0023104, 
    -0.0023104, -0.004501875, -0.005520921, -0.0001224955, 2.964231e-05,
  2.744877e-05, -0.000102832, -0.001694225, -0.0008165565, -0.0001343212, 
    -0.0001343212, -0.0008165565, -0.001694225, -0.000102832, 2.744877e-05,
  -2.744877e-05, 0.000102832, 0.001694225, 0.0008165565, 0.0001343212, 
    0.0001343212, 0.0008165565, 0.001694225, 0.000102832, -2.744877e-05,
  -2.964231e-05, 0.0001224955, 0.005520921, 0.004501875, 0.0023104, 
    0.0023104, 0.004501875, 0.005520921, 0.0001224955, -2.964231e-05,
  0, 0.0002219629, 0.008224508, 0.009216779, 0.009496097, 0.009496097, 
    0.009216779, 0.008224508, 0.0002219629, 0,
  0, 0, 0.0006440201, 0.002197089, 0.00343237, 0.00343237, 0.002197089, 
    0.0006440201, 0, 0,
  0, 0, 0, -0.0005892332, -0.0009190909, -0.0009190909, -0.0005892332, 0, 0, 0,
  0, 0, 0, 0.0005568951, 0.0008832509, 0.0008832509, 0.0005568951, 0, 0, 0,
  0, 0, -0.0005246762, -0.002076827, -0.003296289, -0.003296289, 
    -0.002076827, -0.0005246762, 0, 0,
  0, -0.0001431774, -0.007956518, -0.008900011, -0.009123077, -0.009123077, 
    -0.008900011, -0.007956518, -0.0001431774, 0,
  2.667872e-05, -0.0001096674, -0.005323435, -0.004267382, -0.002119857, 
    -0.002119857, -0.004267382, -0.005323435, -0.0001096674, 2.667872e-05,
  2.664079e-05, -9.966083e-05, -0.001625223, -0.0007479631, -0.0001177278, 
    -0.0001177278, -0.0007479631, -0.001625223, -9.966083e-05, 2.664079e-05,
  -2.664079e-05, 9.966083e-05, 0.001625223, 0.0007479631, 0.0001177278, 
    0.0001177278, 0.0007479631, 0.001625223, 9.966083e-05, -2.664079e-05,
  -2.667872e-05, 0.0001096674, 0.005323435, 0.004267382, 0.002119857, 
    0.002119857, 0.004267382, 0.005323435, 0.0001096674, -2.667872e-05,
  0, 0.0001431774, 0.007956518, 0.008900011, 0.009123077, 0.009123077, 
    0.008900011, 0.007956518, 0.0001431774, 0,
  0, 0, 0.0005246762, 0.002076827, 0.003296289, 0.003296289, 0.002076827, 
    0.0005246762, 0, 0,
  0, 0, 0, -0.0005568951, -0.0008832509, -0.0008832509, -0.0005568951, 0, 0, 0,
  0, 0, 0, 0.0005037647, 0.0008088268, 0.0008088268, 0.0005037647, 0, 0, 0,
  0, 0, -0.0004079585, -0.001878764, -0.00301774, -0.00301774, -0.001878764, 
    -0.0004079585, 0, 0,
  0, -7.64058e-05, -0.007352239, -0.008238082, -0.008422702, -0.008422702, 
    -0.008238082, -0.007352239, -7.64058e-05, 0,
  2.307964e-05, -9.385345e-05, -0.004917953, -0.003885338, -0.001871772, 
    -0.001871772, -0.003885338, -0.004917953, -9.385345e-05, 2.307964e-05,
  2.435831e-05, -9.109949e-05, -0.001498217, -0.00066039, -9.806082e-05, 
    -9.806082e-05, -0.00066039, -0.001498217, -9.109949e-05, 2.435831e-05,
  -2.435831e-05, 9.109949e-05, 0.001498217, 0.00066039, 9.806082e-05, 
    9.806082e-05, 0.00066039, 0.001498217, 9.109949e-05, -2.435831e-05,
  -2.307964e-05, 9.385345e-05, 0.004917953, 0.003885338, 0.001871772, 
    0.001871772, 0.003885338, 0.004917953, 9.385345e-05, -2.307964e-05,
  0, 7.64058e-05, 0.007352239, 0.008238082, 0.008422702, 0.008422702, 
    0.008238082, 0.007352239, 7.64058e-05, 0,
  0, 0, 0.0004079585, 0.001878764, 0.00301774, 0.00301774, 0.001878764, 
    0.0004079585, 0, 0,
  0, 0, 0, -0.0005037647, -0.0008088268, -0.0008088268, -0.0005037647, 0, 0, 0,
  0, 0, 0, 0.0004322374, 0.0006996897, 0.0006996897, 0.0004322374, 0, 0, 0,
  0, 0, -0.0003049664, -0.001612117, -0.002610353, -0.002610353, 
    -0.001612117, -0.0003049664, 0, 0,
  0, -2.918386e-05, -0.006424312, -0.007218394, -0.007378257, -0.007378257, 
    -0.007218394, -0.006424312, -2.918386e-05, 0,
  1.903953e-05, -7.647537e-05, -0.004300881, -0.003362936, -0.001585539, 
    -0.001585539, -0.003362936, -0.004300881, -7.647537e-05, 1.903953e-05,
  2.092772e-05, -7.825991e-05, -0.001310519, -0.0005603368, -7.892161e-05, 
    -7.892161e-05, -0.0005603368, -0.001310519, -7.825991e-05, 2.092772e-05,
  -2.092772e-05, 7.825991e-05, 0.001310519, 0.0005603368, 7.892161e-05, 
    7.892161e-05, 0.0005603368, 0.001310519, 7.825991e-05, -2.092772e-05,
  -1.903953e-05, 7.647537e-05, 0.004300881, 0.003362936, 0.001585539, 
    0.001585539, 0.003362936, 0.004300881, 7.647537e-05, -1.903953e-05,
  0, 2.918386e-05, 0.006424312, 0.007218394, 0.007378257, 0.007378257, 
    0.007218394, 0.006424312, 2.918386e-05, 0,
  0, 0, 0.0003049664, 0.001612117, 0.002610353, 0.002610353, 0.001612117, 
    0.0003049664, 0, 0,
  0, 0, 0, -0.0004322374, -0.0006996897, -0.0006996897, -0.0004322374, 0, 0, 0,
  0, 0, 0, 0.0003490069, 0.0005682205, 0.0005682205, 0.0003490069, 0, 0, 0,
  0, 0, -0.0002173395, -0.001301814, -0.002119897, -0.002119897, 
    -0.001301814, -0.0002173395, 0, 0,
  0, 2.02782e-07, -0.005269258, -0.005936124, -0.00607133, -0.00607133, 
    -0.005936124, -0.005269258, 2.02782e-07, 0,
  1.486524e-05, -5.895624e-05, -0.003530692, -0.002739154, -0.001272735, 
    -0.001272735, -0.002739154, -0.003530692, -5.895624e-05, 1.486524e-05,
  1.686389e-05, -6.30493e-05, -0.00107686, -0.0004509174, -6.133533e-05, 
    -6.133533e-05, -0.0004509174, -0.00107686, -6.30493e-05, 1.686389e-05,
  -1.686389e-05, 6.30493e-05, 0.00107686, 0.0004509174, 6.133533e-05, 
    6.133533e-05, 0.0004509174, 0.00107686, 6.30493e-05, -1.686389e-05,
  -1.486524e-05, 5.895624e-05, 0.003530692, 0.002739154, 0.001272735, 
    0.001272735, 0.002739154, 0.003530692, 5.895624e-05, -1.486524e-05,
  0, -2.02782e-07, 0.005269258, 0.005936124, 0.00607133, 0.00607133, 
    0.005936124, 0.005269258, -2.02782e-07, 0,
  0, 0, 0.0002173395, 0.001301814, 0.002119897, 0.002119897, 0.001301814, 
    0.0002173395, 0, 0,
  0, 0, 0, -0.0003490069, -0.0005682205, -0.0005682205, -0.0003490069, 0, 0, 0,
  0, 0, 0, 0.000260449, 0.0004257144, 0.0004257144, 0.000260449, 0, 0, 0,
  0, 0, -0.0001452263, -0.0009715913, -0.001588321, -0.001588321, 
    -0.0009715913, -0.0001452263, 0, 0,
  0, 1.449837e-05, -0.003986346, -0.004500266, -0.004606354, -0.004606354, 
    -0.004500266, -0.003986346, 1.449837e-05, 0,
  1.078954e-05, -4.224362e-05, -0.00267257, -0.00205993, -0.0009472928, 
    -0.0009472928, -0.00205993, -0.00267257, -4.224362e-05, 1.078954e-05,
  1.253975e-05, -4.68675e-05, -0.0008159337, -0.0003365328, -4.491138e-05, 
    -4.491138e-05, -0.0003365328, -0.0008159337, -4.68675e-05, 1.253975e-05,
  -1.253975e-05, 4.68675e-05, 0.0008159337, 0.0003365328, 4.491138e-05, 
    4.491138e-05, 0.0003365328, 0.0008159337, 4.68675e-05, -1.253975e-05,
  -1.078954e-05, 4.224362e-05, 0.00267257, 0.00205993, 0.0009472928, 
    0.0009472928, 0.00205993, 0.00267257, 4.224362e-05, -1.078954e-05,
  0, -1.449837e-05, 0.003986346, 0.004500266, 0.004606354, 0.004606354, 
    0.004500266, 0.003986346, -1.449837e-05, 0,
  0, 0, 0.0001452263, 0.0009715913, 0.001588321, 0.001588321, 0.0009715913, 
    0.0001452263, 0, 0,
  0, 0, 0, -0.000260449, -0.0004257144, -0.0004257144, -0.000260449, 0, 0, 0,
  0, 0, 0, 0.0001711433, 0.0002804244, 0.0002804244, 0.0001711433, 0, 0, 0,
  0, 0, -8.680863e-05, -0.0006385141, -0.001046328, -0.001046328, 
    -0.0006385141, -8.680863e-05, 0, 0,
  0, 1.717206e-05, -0.002652172, -0.002999044, -0.003071944, -0.003071944, 
    -0.002999044, -0.002652172, 1.717206e-05, 0,
  6.926054e-06, -2.675768e-05, -0.001778646, -0.001362896, -0.0006218205, 
    -0.0006218205, -0.001362896, -0.001778646, -2.675768e-05, 6.926054e-06,
  8.20167e-06, -3.064086e-05, -0.0005434534, -0.0002215119, -2.930621e-05, 
    -2.930621e-05, -0.0002215119, -0.0005434534, -3.064086e-05, 8.20167e-06,
  -8.20167e-06, 3.064086e-05, 0.0005434534, 0.0002215119, 2.930621e-05, 
    2.930621e-05, 0.0002215119, 0.0005434534, 3.064086e-05, -8.20167e-06,
  -6.926054e-06, 2.675768e-05, 0.001778646, 0.001362896, 0.0006218205, 
    0.0006218205, 0.001362896, 0.001778646, 2.675768e-05, -6.926054e-06,
  0, -1.717206e-05, 0.002652172, 0.002999044, 0.003071944, 0.003071944, 
    0.002999044, 0.002652172, -1.717206e-05, 0,
  0, 0, 8.680863e-05, 0.0006385141, 0.001046328, 0.001046328, 0.0006385141, 
    8.680863e-05, 0, 0,
  0, 0, 0, -0.0001711433, -0.0002804244, -0.0002804244, -0.0001711433, 0, 0, 0,
  0, 0, 0, 8.384304e-05, 0.0001376203, 0.0001376203, 8.384304e-05, 0, 0, 0,
  0, 0, -3.896345e-05, -0.0003128497, -0.0005135435, -0.0005135435, 
    -0.0003128497, -3.896345e-05, 0, 0,
  0, 1.176195e-05, -0.001315608, -0.001491015, -0.001528998, -0.001528998, 
    -0.001491015, -0.001315608, 1.176195e-05, 0,
  3.30618e-06, -1.258667e-05, -0.0008832358, -0.000673676, -0.0003052508, 
    -0.0003052508, -0.000673676, -0.0008832358, -1.258667e-05, 3.30618e-06,
  3.997906e-06, -1.492714e-05, -0.0002701678, -0.0001090037, -1.43951e-05, 
    -1.43951e-05, -0.0001090037, -0.0002701678, -1.492714e-05, 3.997906e-06,
  -3.997906e-06, 1.492714e-05, 0.0002701678, 0.0001090037, 1.43951e-05, 
    1.43951e-05, 0.0001090037, 0.0002701678, 1.492714e-05, -3.997906e-06,
  -3.30618e-06, 1.258667e-05, 0.0008832358, 0.000673676, 0.0003052508, 
    0.0003052508, 0.000673676, 0.0008832358, 1.258667e-05, -3.30618e-06,
  0, -1.176195e-05, 0.001315608, 0.001491015, 0.001528998, 0.001528998, 
    0.001491015, 0.001315608, -1.176195e-05, 0,
  0, 0, 3.896345e-05, 0.0003128497, 0.0005135435, 0.0005135435, 0.0003128497, 
    3.896345e-05, 0, 0,
  0, 0, 0, -8.384304e-05, -0.0001376203, -0.0001376203, -8.384304e-05, 0, 0, 0,
  0, 0, 0, 5.815344e-09, 7.002647e-09, 7.002647e-09, 5.815344e-09, 0, 0, 0,
  0, 0, -1.32585e-08, -2.381267e-08, -2.868336e-08, -2.868336e-08, 
    -2.381267e-08, -1.32585e-08, 0, 0,
  0, -1.15415e-08, -2.346004e-08, -2.459297e-08, -2.537498e-08, 
    -2.537498e-08, -2.459297e-08, -2.346004e-08, -1.15415e-08, 0,
  5.857667e-10, -4.246539e-09, -1.556134e-08, -1.540685e-08, -1.532166e-08, 
    -1.532166e-08, -1.540685e-08, -1.556134e-08, -4.246539e-09, 5.857667e-10,
  3.120892e-10, -1.097673e-09, -4.869617e-09, -5.098232e-09, -5.842038e-09, 
    -5.842038e-09, -5.098232e-09, -4.869617e-09, -1.097673e-09, 3.120892e-10,
  -3.120892e-10, 1.097673e-09, 4.869617e-09, 5.098232e-09, 5.842038e-09, 
    5.842038e-09, 5.098232e-09, 4.869617e-09, 1.097673e-09, -3.120892e-10,
  -5.857667e-10, 4.246539e-09, 1.556134e-08, 1.540685e-08, 1.532166e-08, 
    1.532166e-08, 1.540685e-08, 1.556134e-08, 4.246539e-09, -5.857667e-10,
  0, 1.15415e-08, 2.346004e-08, 2.459297e-08, 2.537498e-08, 2.537498e-08, 
    2.459297e-08, 2.346004e-08, 1.15415e-08, 0,
  0, 0, 1.32585e-08, 2.381267e-08, 2.868336e-08, 2.868336e-08, 2.381267e-08, 
    1.32585e-08, 0, 0,
  0, 0, 0, -5.815344e-09, -7.002647e-09, -7.002647e-09, -5.815344e-09, 0, 0, 0,
  0, 0, 0, 0.0006061294, 0.0009345636, 0.0009345636, 0.0006061294, 0, 0, 0,
  0, 0, -0.00072758, -0.002260444, -0.00349472, -0.00349472, -0.002260444, 
    -0.00072758, 0, 0,
  0, -0.0002768362, -0.008301422, -0.009286314, -0.009566539, -0.009566539, 
    -0.009286314, -0.008301422, -0.0002768362, 0,
  3.247311e-05, -0.0001333559, -0.005568251, -0.004563344, -0.002390856, 
    -0.002390856, -0.004563344, -0.005568251, -0.0001333559, 3.247311e-05,
  2.790047e-05, -0.0001046175, -0.001709754, -0.0008484946, -0.000145277, 
    -0.000145277, -0.0008484946, -0.001709754, -0.0001046175, 2.790047e-05,
  -2.790047e-05, 0.0001046175, 0.001709754, 0.0008484946, 0.000145277, 
    0.000145277, 0.0008484946, 0.001709754, 0.0001046175, -2.790047e-05,
  -3.247311e-05, 0.0001333559, 0.005568251, 0.004563344, 0.002390856, 
    0.002390856, 0.004563344, 0.005568251, 0.0001333559, -3.247311e-05,
  0, 0.0002768362, 0.008301422, 0.009286314, 0.009566539, 0.009566539, 
    0.009286314, 0.008301422, 0.0002768362, 0,
  0, 0, 0.00072758, 0.002260444, 0.00349472, 0.00349472, 0.002260444, 
    0.00072758, 0, 0,
  0, 0, 0, -0.0006061294, -0.0009345636, -0.0009345636, -0.0006061294, 0, 0, 0,
  0, 0, 0, 0.0005934635, 0.000923071, 0.000923071, 0.0005934635, 0, 0, 0,
  0, 0, -0.0006609037, -0.002212907, -0.003447313, -0.003447313, 
    -0.002212907, -0.0006609037, 0, 0,
  0, -0.0002331512, -0.008230937, -0.009184726, -0.009438962, -0.009438962, 
    -0.009184726, -0.008230937, -0.0002331512, 0,
  3.064858e-05, -0.0001262809, -0.005506466, -0.004486478, -0.002315367, 
    -0.002315367, -0.004486478, -0.005506466, -0.0001262809, 3.064858e-05,
  2.766737e-05, -0.0001036354, -0.001686466, -0.0008188451, -0.0001367709, 
    -0.0001367709, -0.0008188451, -0.001686466, -0.0001036354, 2.766737e-05,
  -2.766737e-05, 0.0001036354, 0.001686466, 0.0008188451, 0.0001367709, 
    0.0001367709, 0.0008188451, 0.001686466, 0.0001036354, -2.766737e-05,
  -3.064858e-05, 0.0001262809, 0.005506466, 0.004486478, 0.002315367, 
    0.002315367, 0.004486478, 0.005506466, 0.0001262809, -3.064858e-05,
  0, 0.0002331512, 0.008230937, 0.009184726, 0.009438962, 0.009438962, 
    0.009184726, 0.008230937, 0.0002331512, 0,
  0, 0, 0.0006609037, 0.002212907, 0.003447313, 0.003447313, 0.002212907, 
    0.0006609037, 0, 0,
  0, 0, 0, -0.0005934635, -0.000923071, -0.000923071, -0.0005934635, 0, 0, 0,
  0, 0, 0, 0.0005610802, 0.0008871742, 0.0008871742, 0.0005610802, 0, 0, 0,
  0, 0, -0.0005412701, -0.002092445, -0.003310974, -0.003310974, 
    -0.002092445, -0.0005412701, 0, 0,
  0, -0.0001542188, -0.007963161, -0.008869411, -0.009069029, -0.009069029, 
    -0.008869411, -0.007963161, -0.0001542188, 0,
  2.767257e-05, -0.0001133935, -0.005309715, -0.004252854, -0.002125125, 
    -0.002125125, -0.004252854, -0.005309715, -0.0001133935, 2.767257e-05,
  2.685105e-05, -0.0001004356, -0.001617949, -0.0007504071, -0.0001198822, 
    -0.0001198822, -0.0007504071, -0.001617949, -0.0001004356, 2.685105e-05,
  -2.685105e-05, 0.0001004356, 0.001617949, 0.0007504071, 0.0001198822, 
    0.0001198822, 0.0007504071, 0.001617949, 0.0001004356, -2.685105e-05,
  -2.767257e-05, 0.0001133935, 0.005309715, 0.004252854, 0.002125125, 
    0.002125125, 0.004252854, 0.005309715, 0.0001133935, -2.767257e-05,
  0, 0.0001542188, 0.007963161, 0.008869411, 0.009069029, 0.009069029, 
    0.008869411, 0.007963161, 0.0001542188, 0,
  0, 0, 0.0005412701, 0.002092445, 0.003310974, 0.003310974, 0.002092445, 
    0.0005412701, 0, 0,
  0, 0, 0, -0.0005610802, -0.0008871742, -0.0008871742, -0.0005610802, 0, 0, 0,
  0, 0, 0, 0.000507704, 0.0008125075, 0.0008125075, 0.000507704, 0, 0, 0,
  0, 0, -0.0004234944, -0.001893454, -0.003031498, -0.003031498, 
    -0.001893454, -0.0004234944, 0, 0,
  0, -8.674272e-05, -0.007359335, -0.008210418, -0.008373619, -0.008373619, 
    -0.008210418, -0.007359335, -8.674272e-05, 0,
  2.400551e-05, -9.731921e-05, -0.004905664, -0.003872271, -0.001877165, 
    -0.001877165, -0.003872271, -0.004905664, -9.731921e-05, 2.400551e-05,
  2.455148e-05, -9.181334e-05, -0.001491658, -0.0006628838, -9.98738e-05, 
    -9.98738e-05, -0.0006628838, -0.001491658, -9.181334e-05, 2.455148e-05,
  -2.455148e-05, 9.181334e-05, 0.001491658, 0.0006628838, 9.98738e-05, 
    9.98738e-05, 0.0006628838, 0.001491658, 9.181334e-05, -2.455148e-05,
  -2.400551e-05, 9.731921e-05, 0.004905664, 0.003872271, 0.001877165, 
    0.001877165, 0.003872271, 0.004905664, 9.731921e-05, -2.400551e-05,
  0, 8.674272e-05, 0.007359335, 0.008210418, 0.008373619, 0.008373619, 
    0.008210418, 0.007359335, 8.674272e-05, 0,
  0, 0, 0.0004234944, 0.001893454, 0.003031498, 0.003031498, 0.001893454, 
    0.0004234944, 0, 0,
  0, 0, 0, -0.000507704, -0.0008125075, -0.0008125075, -0.000507704, 0, 0, 0,
  0, 0, 0, 0.0004357429, 0.0007029631, 0.0007029631, 0.0004357429, 0, 0, 0,
  0, 0, -0.0003187215, -0.001625186, -0.002622579, -0.002622579, 
    -0.001625186, -0.0003187215, 0, 0,
  0, -3.829163e-05, -0.006431939, -0.007195233, -0.007336242, -0.007336242, 
    -0.007195233, -0.006431939, -3.829163e-05, 0,
  1.984986e-05, -7.950608e-05, -0.004290752, -0.003351852, -0.001590661, 
    -0.001590661, -0.003351852, -0.004290752, -7.950608e-05, 1.984986e-05,
  2.109633e-05, -7.888443e-05, -0.001304943, -0.000562699, -8.040916e-05, 
    -8.040916e-05, -0.000562699, -0.001304943, -7.888443e-05, 2.109633e-05,
  -2.109633e-05, 7.888443e-05, 0.001304943, 0.000562699, 8.040916e-05, 
    8.040916e-05, 0.000562699, 0.001304943, 7.888443e-05, -2.109633e-05,
  -1.984986e-05, 7.950608e-05, 0.004290752, 0.003351852, 0.001590661, 
    0.001590661, 0.003351852, 0.004290752, 7.950608e-05, -1.984986e-05,
  0, 3.829163e-05, 0.006431939, 0.007195233, 0.007336242, 0.007336242, 
    0.007195233, 0.006431939, 3.829163e-05, 0,
  0, 0, 0.0003187215, 0.001625186, 0.002622579, 0.002622579, 0.001625186, 
    0.0003187215, 0, 0,
  0, 0, 0, -0.0004357429, -0.0007029631, -0.0007029631, -0.0004357429, 0, 0, 0,
  0, 0, 0, 0.0003519526, 0.000570968, 0.000570968, 0.0003519526, 0, 0, 0,
  0, 0, -0.0002288451, -0.001312796, -0.002130154, -0.002130154, 
    -0.001312796, -0.0002288451, 0, 0,
  0, -7.34213e-06, -0.005277331, -0.005918587, -0.006038046, -0.006038046, 
    -0.005918587, -0.005277331, -7.34213e-06, 0,
  1.552998e-05, -6.144099e-05, -0.003523243, -0.00273045, -0.001277258, 
    -0.001277258, -0.00273045, -0.003523243, -6.144099e-05, 1.552998e-05,
  1.700224e-05, -6.356273e-05, -0.001072489, -0.0004529995, -6.251538e-05, 
    -6.251538e-05, -0.0004529995, -0.001072489, -6.356273e-05, 1.700224e-05,
  -1.700224e-05, 6.356273e-05, 0.001072489, 0.0004529995, 6.251538e-05, 
    6.251538e-05, 0.0004529995, 0.001072489, 6.356273e-05, -1.700224e-05,
  -1.552998e-05, 6.144099e-05, 0.003523243, 0.00273045, 0.001277258, 
    0.001277258, 0.00273045, 0.003523243, 6.144099e-05, -1.552998e-05,
  0, 7.34213e-06, 0.005277331, 0.005918587, 0.006038046, 0.006038046, 
    0.005918587, 0.005277331, 7.34213e-06, 0,
  0, 0, 0.0002288451, 0.001312796, 0.002130154, 0.002130154, 0.001312796, 
    0.0002288451, 0, 0,
  0, 0, 0, -0.0003519526, -0.000570968, -0.000570968, -0.0003519526, 0, 0, 0,
  0, 0, 0, 0.0002627548, 0.0004278635, 0.0004278635, 0.0002627548, 0, 0, 0,
  0, 0, -0.0001541701, -0.0009801878, -0.001596342, -0.001596342, 
    -0.0009801878, -0.0001541701, 0, 0,
  0, 8.722372e-06, -0.003994514, -0.004488886, -0.004582806, -0.004582806, 
    -0.004488886, -0.003994514, 8.722372e-06, 0,
  1.129161e-05, -4.411942e-05, -0.002668035, -0.002053865, -0.0009510084, 
    -0.0009510084, -0.002053865, -0.002668035, -4.411942e-05, 1.129161e-05,
  1.264471e-05, -4.725766e-05, -0.0008129022, -0.0003382375, -4.579626e-05, 
    -4.579626e-05, -0.0003382375, -0.0008129022, -4.725766e-05, 1.264471e-05,
  -1.264471e-05, 4.725766e-05, 0.0008129022, 0.0003382375, 4.579626e-05, 
    4.579626e-05, 0.0003382375, 0.0008129022, 4.725766e-05, -1.264471e-05,
  -1.129161e-05, 4.411942e-05, 0.002668035, 0.002053865, 0.0009510084, 
    0.0009510084, 0.002053865, 0.002668035, 4.411942e-05, -1.129161e-05,
  0, -8.722372e-06, 0.003994514, 0.004488886, 0.004582806, 0.004582806, 
    0.004488886, 0.003994514, -8.722372e-06, 0,
  0, 0, 0.0001541701, 0.0009801878, 0.001596342, 0.001596342, 0.0009801878, 
    0.0001541701, 0, 0,
  0, 0, 0, -0.0002627548, -0.0004278635, -0.0004278635, -0.0002627548, 0, 0, 0,
  0, 0, 0, 0.0001727396, 0.0002819296, 0.0002819296, 0.0001727396, 0, 0, 0,
  0, 0, -9.286299e-05, -0.0006444664, -0.001051945, -0.001051945, 
    -0.0006444664, -9.286299e-05, 0, 0,
  0, 1.334456e-05, -0.002659449, -0.002993557, -0.003058342, -0.003058342, 
    -0.002993557, -0.002659449, 1.334456e-05, 0,
  7.255041e-06, -2.798641e-05, -0.001776851, -0.001359622, -0.0006246124, 
    -0.0006246124, -0.001359622, -0.001776851, -2.798641e-05, 7.255041e-06,
  8.272434e-06, -3.090431e-05, -0.0005417906, -0.000222772, -2.990525e-05, 
    -2.990525e-05, -0.000222772, -0.0005417906, -3.090431e-05, 8.272434e-06,
  -8.272434e-06, 3.090431e-05, 0.0005417906, 0.000222772, 2.990525e-05, 
    2.990525e-05, 0.000222772, 0.0005417906, 3.090431e-05, -8.272434e-06,
  -7.255041e-06, 2.798641e-05, 0.001776851, 0.001359622, 0.0006246124, 
    0.0006246124, 0.001359622, 0.001776851, 2.798641e-05, -7.255041e-06,
  0, -1.334456e-05, 0.002659449, 0.002993557, 0.003058342, 0.003058342, 
    0.002993557, 0.002659449, -1.334456e-05, 0,
  0, 0, 9.286299e-05, 0.0006444664, 0.001051945, 0.001051945, 0.0006444664, 
    9.286299e-05, 0, 0,
  0, 0, 0, -0.0001727396, -0.0002819296, -0.0002819296, -0.0001727396, 0, 0, 0,
  0, 0, 0, 8.465277e-05, 0.000138414, 0.000138414, 8.465277e-05, 0, 0, 0,
  0, 0, -4.188015e-05, -0.0003158701, -0.0005165051, -0.0005165051, 
    -0.0003158701, -4.188015e-05, 0, 0,
  0, 9.967926e-06, -0.00132016, -0.001489761, -0.001523985, -0.001523985, 
    -0.001489761, -0.00132016, 9.967926e-06, 0,
  3.460302e-06, -1.316213e-05, -0.0008832128, -0.000672873, -0.0003069691, 
    -0.0003069691, -0.000672873, -0.0008832128, -1.316213e-05, 3.460302e-06,
  4.033622e-06, -1.50603e-05, -0.0002696476, -0.0001097427, -1.470675e-05, 
    -1.470675e-05, -0.0001097427, -0.0002696476, -1.50603e-05, 4.033622e-06,
  -4.033622e-06, 1.50603e-05, 0.0002696476, 0.0001097427, 1.470675e-05, 
    1.470675e-05, 0.0001097427, 0.0002696476, 1.50603e-05, -4.033622e-06,
  -3.460302e-06, 1.316213e-05, 0.0008832128, 0.000672873, 0.0003069691, 
    0.0003069691, 0.000672873, 0.0008832128, 1.316213e-05, -3.460302e-06,
  0, -9.967926e-06, 0.00132016, 0.001489761, 0.001523985, 0.001523985, 
    0.001489761, 0.00132016, -9.967926e-06, 0,
  0, 0, 4.188015e-05, 0.0003158701, 0.0005165051, 0.0005165051, 0.0003158701, 
    4.188015e-05, 0, 0,
  0, 0, 0, -8.465277e-05, -0.000138414, -0.000138414, -8.465277e-05, 0, 0, 0,
  0, 0, 0, 5.818711e-09, 7.003219e-09, 7.003219e-09, 5.818711e-09, 0, 0, 0,
  0, 0, -1.328672e-08, -2.384211e-08, -2.870693e-08, -2.870693e-08, 
    -2.384211e-08, -1.328672e-08, 0, 0,
  0, -1.155473e-08, -2.345341e-08, -2.454256e-08, -2.530428e-08, 
    -2.530428e-08, -2.454256e-08, -2.345341e-08, -1.155473e-08, 0,
  5.859639e-10, -4.252366e-09, -1.554851e-08, -1.538936e-08, -1.532886e-08, 
    -1.532886e-08, -1.538936e-08, -1.554851e-08, -4.252366e-09, 5.859639e-10,
  3.12195e-10, -1.098231e-09, -4.866877e-09, -5.100642e-09, -5.862804e-09, 
    -5.862804e-09, -5.100642e-09, -4.866877e-09, -1.098231e-09, 3.12195e-10,
  -3.12195e-10, 1.098231e-09, 4.866877e-09, 5.100642e-09, 5.862804e-09, 
    5.862804e-09, 5.100642e-09, 4.866877e-09, 1.098231e-09, -3.12195e-10,
  -5.859639e-10, 4.252366e-09, 1.554851e-08, 1.538936e-08, 1.532886e-08, 
    1.532886e-08, 1.538936e-08, 1.554851e-08, 4.252366e-09, -5.859639e-10,
  0, 1.155473e-08, 2.345341e-08, 2.454256e-08, 2.530428e-08, 2.530428e-08, 
    2.454256e-08, 2.345341e-08, 1.155473e-08, 0,
  0, 0, 1.328672e-08, 2.384211e-08, 2.870693e-08, 2.870693e-08, 2.384211e-08, 
    1.328672e-08, 0, 0,
  0, 0, 0, -5.818711e-09, -7.003219e-09, -7.003219e-09, -5.818711e-09, 0, 0, 0,
  0, 0, 0, 0.0006103343, 0.0009384871, 0.0009384871, 0.0006103343, 0, 0, 0,
  0, 0, -0.0007443273, -0.002276226, -0.003509531, -0.003509531, 
    -0.002276226, -0.0007443273, 0, 0,
  0, -0.0002879208, -0.008307651, -0.00925385, -0.009508641, -0.009508641, 
    -0.00925385, -0.008307651, -0.0002879208, 0,
  3.347251e-05, -0.0001371278, -0.005553571, -0.004547864, -0.002395635, 
    -0.002395635, -0.004547864, -0.005553571, -0.0001371278, 3.347251e-05,
  2.81193e-05, -0.0001054216, -0.001701849, -0.0008506518, -0.0001478502, 
    -0.0001478502, -0.0008506518, -0.001701849, -0.0001054216, 2.81193e-05,
  -2.81193e-05, 0.0001054216, 0.001701849, 0.0008506518, 0.0001478502, 
    0.0001478502, 0.0008506518, 0.001701849, 0.0001054216, -2.81193e-05,
  -3.347251e-05, 0.0001371278, 0.005553571, 0.004547864, 0.002395635, 
    0.002395635, 0.004547864, 0.005553571, 0.0001371278, -3.347251e-05,
  0, 0.0002879208, 0.008307651, 0.00925385, 0.009508641, 0.009508641, 
    0.00925385, 0.008307651, 0.0002879208, 0,
  0, 0, 0.0007443273, 0.002276226, 0.003509531, 0.003509531, 0.002276226, 
    0.0007443273, 0, 0,
  0, 0, 0, -0.0006103343, -0.0009384871, -0.0009384871, -0.0006103343, 0, 0, 0,
  0, 0, 0, 0.0005976752, 0.0009270158, 0.0009270158, 0.0005976752, 0, 0, 0,
  0, 0, -0.0006777684, -0.002228657, -0.003462126, -0.003462126, 
    -0.002228657, -0.0006777684, 0, 0,
  0, -0.0002443254, -0.008237146, -0.009152789, -0.00938243, -0.00938243, 
    -0.009152789, -0.008237146, -0.0002443254, 0,
  3.165267e-05, -0.000130058, -0.00549205, -0.004471213, -0.002320217, 
    -0.002320217, -0.004471213, -0.00549205, -0.000130058, 3.165267e-05,
  2.788437e-05, -0.0001044329, -0.001678783, -0.000821099, -0.0001392249, 
    -0.0001392249, -0.000821099, -0.001678783, -0.0001044329, 2.788437e-05,
  -2.788437e-05, 0.0001044329, 0.001678783, 0.000821099, 0.0001392249, 
    0.0001392249, 0.000821099, 0.001678783, 0.0001044329, -2.788437e-05,
  -3.165267e-05, 0.000130058, 0.00549205, 0.004471213, 0.002320217, 
    0.002320217, 0.004471213, 0.00549205, 0.000130058, -3.165267e-05,
  0, 0.0002443254, 0.008237146, 0.009152789, 0.00938243, 0.00938243, 
    0.009152789, 0.008237146, 0.0002443254, 0,
  0, 0, 0.0006777684, 0.002228657, 0.003462126, 0.003462126, 0.002228657, 
    0.0006777684, 0, 0,
  0, 0, 0, -0.0005976752, -0.0009270158, -0.0009270158, -0.0005976752, 0, 0, 0,
  0, 0, 0, 0.0005652474, 0.000891063, 0.000891063, 0.0005652474, 0, 0, 0,
  0, 0, -0.0005578496, -0.002107996, -0.003325532, -0.003325532, 
    -0.002107996, -0.0005578496, 0, 0,
  0, -0.0001652497, -0.007969586, -0.008838919, -0.009015546, -0.009015546, 
    -0.008838919, -0.007969586, -0.0001652497, 0,
  2.866435e-05, -0.0001171117, -0.005296031, -0.004238452, -0.00213028, 
    -0.00213028, -0.004238452, -0.005296031, -0.0001171117, 2.866435e-05,
  2.705974e-05, -0.0001012046, -0.001610746, -0.0007528162, -0.0001220418, 
    -0.0001220418, -0.0007528162, -0.001610746, -0.0001012046, 2.705974e-05,
  -2.705974e-05, 0.0001012046, 0.001610746, 0.0007528162, 0.0001220418, 
    0.0001220418, 0.0007528162, 0.001610746, 0.0001012046, -2.705974e-05,
  -2.866435e-05, 0.0001171117, 0.005296031, 0.004238452, 0.00213028, 
    0.00213028, 0.004238452, 0.005296031, 0.0001171117, -2.866435e-05,
  0, 0.0001652497, 0.007969586, 0.008838919, 0.009015546, 0.009015546, 
    0.008838919, 0.007969586, 0.0001652497, 0,
  0, 0, 0.0005578496, 0.002107996, 0.003325532, 0.003325532, 0.002107996, 
    0.0005578496, 0, 0,
  0, 0, 0, -0.0005652474, -0.000891063, -0.000891063, -0.0005652474, 0, 0, 0,
  0, 0, 0, 0.0005116269, 0.0008161564, 0.0008161564, 0.0005116269, 0, 0, 0,
  0, 0, -0.0004390201, -0.001908083, -0.003045139, -0.003045139, 
    -0.001908083, -0.0004390201, 0, 0,
  0, -9.707255e-05, -0.007366215, -0.00818284, -0.008325042, -0.008325042, 
    -0.00818284, -0.007366215, -9.707255e-05, 0,
  2.492957e-05, -0.000100778, -0.004893403, -0.003859318, -0.001882452, 
    -0.001882452, -0.003859318, -0.004893403, -0.000100778, 2.492957e-05,
  2.474323e-05, -9.252194e-05, -0.001485162, -0.0006653439, -0.0001016929, 
    -0.0001016929, -0.0006653439, -0.001485162, -9.252194e-05, 2.474323e-05,
  -2.474323e-05, 9.252194e-05, 0.001485162, 0.0006653439, 0.0001016929, 
    0.0001016929, 0.0006653439, 0.001485162, 9.252194e-05, -2.474323e-05,
  -2.492957e-05, 0.000100778, 0.004893403, 0.003859318, 0.001882452, 
    0.001882452, 0.003859318, 0.004893403, 0.000100778, -2.492957e-05,
  0, 9.707255e-05, 0.007366215, 0.00818284, 0.008325042, 0.008325042, 
    0.00818284, 0.007366215, 9.707255e-05, 0,
  0, 0, 0.0004390201, 0.001908083, 0.003045139, 0.003045139, 0.001908083, 
    0.0004390201, 0, 0,
  0, 0, 0, -0.0005116269, -0.0008161564, -0.0008161564, -0.0005116269, 0, 0, 0,
  0, 0, 0, 0.0004392341, 0.0007062089, 0.0007062089, 0.0004392341, 0, 0, 0,
  0, 0, -0.00033247, -0.001638202, -0.002634703, -0.002634703, -0.001638202, 
    -0.00033247, 0, 0,
  0, -4.739587e-05, -0.006439356, -0.007172128, -0.007294649, -0.007294649, 
    -0.007172128, -0.006439356, -4.739587e-05, 0,
  2.065873e-05, -8.253117e-05, -0.004280637, -0.003340868, -0.001595689, 
    -0.001595689, -0.003340868, -0.004280637, -8.253117e-05, 2.065873e-05,
  2.126374e-05, -7.950452e-05, -0.001299421, -0.0005650306, -8.190312e-05, 
    -8.190312e-05, -0.0005650306, -0.001299421, -7.950452e-05, 2.126374e-05,
  -2.126374e-05, 7.950452e-05, 0.001299421, 0.0005650306, 8.190312e-05, 
    8.190312e-05, 0.0005650306, 0.001299421, 7.950452e-05, -2.126374e-05,
  -2.065873e-05, 8.253117e-05, 0.004280637, 0.003340868, 0.001595689, 
    0.001595689, 0.003340868, 0.004280637, 8.253117e-05, -2.065873e-05,
  0, 4.739587e-05, 0.006439356, 0.007172128, 0.007294649, 0.007294649, 
    0.007172128, 0.006439356, 4.739587e-05, 0,
  0, 0, 0.00033247, 0.001638202, 0.002634703, 0.002634703, 0.001638202, 
    0.00033247, 0, 0,
  0, 0, 0, -0.0004392341, -0.0007062089, -0.0007062089, -0.0004392341, 0, 0, 0,
  0, 0, 0, 0.000354886, 0.0005736933, 0.0005736933, 0.000354886, 0, 0, 0,
  0, 0, -0.0002403419, -0.001323731, -0.002140329, -0.002140329, 
    -0.001323731, -0.0002403419, 0, 0,
  0, -1.488402e-05, -0.00528519, -0.005901063, -0.006005088, -0.006005088, 
    -0.005901063, -0.00528519, -1.488402e-05, 0,
  1.619353e-05, -6.392113e-05, -0.003515788, -0.002721828, -0.001281703, 
    -0.001281703, -0.002721828, -0.003515788, -6.392113e-05, 1.619353e-05,
  1.713968e-05, -6.40728e-05, -0.001068158, -0.0004550555, -6.370142e-05, 
    -6.370142e-05, -0.0004550555, -0.001068158, -6.40728e-05, 1.713968e-05,
  -1.713968e-05, 6.40728e-05, 0.001068158, 0.0004550555, 6.370142e-05, 
    6.370142e-05, 0.0004550555, 0.001068158, 6.40728e-05, -1.713968e-05,
  -1.619353e-05, 6.392113e-05, 0.003515788, 0.002721828, 0.001281703, 
    0.001281703, 0.002721828, 0.003515788, 6.392113e-05, -1.619353e-05,
  0, 1.488402e-05, 0.00528519, 0.005901063, 0.006005088, 0.006005088, 
    0.005901063, 0.00528519, 1.488402e-05, 0,
  0, 0, 0.0002403419, 0.001323731, 0.002140329, 0.002140329, 0.001323731, 
    0.0002403419, 0, 0,
  0, 0, 0, -0.000354886, -0.0005736933, -0.0005736933, -0.000354886, 0, 0, 0,
  0, 0, 0, 0.0002650476, 0.0004299959, 0.0004299959, 0.0002650476, 0, 0, 0,
  0, 0, -0.0001630833, -0.0009887358, -0.0016043, -0.0016043, -0.0009887358, 
    -0.0001630833, 0, 0,
  0, 2.959485e-06, -0.004002416, -0.004477448, -0.004559465, -0.004559465, 
    -0.004477448, -0.004002416, 2.959485e-06, 0,
  1.179233e-05, -4.599014e-05, -0.002663461, -0.002047871, -0.0009546667, 
    -0.0009546667, -0.002047871, -0.002663461, -4.599014e-05, 1.179233e-05,
  1.274914e-05, -4.764587e-05, -0.0008098975, -0.0003399205, -4.66862e-05, 
    -4.66862e-05, -0.0003399205, -0.0008098975, -4.764587e-05, 1.274914e-05,
  -1.274914e-05, 4.764587e-05, 0.0008098975, 0.0003399205, 4.66862e-05, 
    4.66862e-05, 0.0003399205, 0.0008098975, 4.764587e-05, -1.274914e-05,
  -1.179233e-05, 4.599014e-05, 0.002663461, 0.002047871, 0.0009546667, 
    0.0009546667, 0.002047871, 0.002663461, 4.599014e-05, -1.179233e-05,
  0, -2.959485e-06, 0.004002416, 0.004477448, 0.004559465, 0.004559465, 
    0.004477448, 0.004002416, -2.959485e-06, 0,
  0, 0, 0.0001630833, 0.0009887358, 0.0016043, 0.0016043, 0.0009887358, 
    0.0001630833, 0, 0,
  0, 0, 0, -0.0002650476, -0.0004299959, -0.0004299959, -0.0002650476, 0, 0, 0,
  0, 0, 0, 0.0001743191, 0.0002834205, 0.0002834205, 0.0001743191, 0, 0, 0,
  0, 0, -9.885567e-05, -0.0006503563, -0.001057508, -0.001057508, 
    -0.0006503563, -9.885567e-05, 0, 0,
  0, 9.544734e-06, -0.002666362, -0.00298789, -0.003044778, -0.003044778, 
    -0.00298789, -0.002666362, 9.544734e-06, 0,
  7.582334e-06, -2.920879e-05, -0.001774951, -0.001356395, -0.0006273668, 
    -0.0006273668, -0.001356395, -0.001774951, -2.920879e-05, 7.582334e-06,
  8.342955e-06, -3.116686e-05, -0.0005401318, -0.0002240145, -3.050758e-05, 
    -3.050758e-05, -0.0002240145, -0.0005401318, -3.116686e-05, 8.342955e-06,
  -8.342955e-06, 3.116686e-05, 0.0005401318, 0.0002240145, 3.050758e-05, 
    3.050758e-05, 0.0002240145, 0.0005401318, 3.116686e-05, -8.342955e-06,
  -7.582334e-06, 2.920879e-05, 0.001774951, 0.001356395, 0.0006273668, 
    0.0006273668, 0.001356395, 0.001774951, 2.920879e-05, -7.582334e-06,
  0, -9.544734e-06, 0.002666362, 0.00298789, 0.003044778, 0.003044778, 
    0.00298789, 0.002666362, -9.544734e-06, 0,
  0, 0, 9.885567e-05, 0.0006503563, 0.001057508, 0.001057508, 0.0006503563, 
    9.885567e-05, 0, 0,
  0, 0, 0, -0.0001743191, -0.0002834205, -0.0002834205, -0.0001743191, 0, 0, 0,
  0, 0, 0, 8.544845e-05, 0.0001391938, 0.0001391938, 8.544845e-05, 0, 0, 0,
  0, 0, -4.47583e-05, -0.0003188381, -0.0005194148, -0.0005194148, 
    -0.0003188381, -4.47583e-05, 0, 0,
  0, 8.185861e-06, -0.001324375, -0.001488222, -0.001518787, -0.001518787, 
    -0.001488222, -0.001324375, 8.185861e-06, 0,
  3.613859e-06, -1.373546e-05, -0.000883024, -0.0006720317, -0.0003086543, 
    -0.0003086543, -0.0006720317, -0.000883024, -1.373546e-05, 3.613859e-06,
  4.069061e-06, -1.519242e-05, -0.0002690957, -0.0001104672, -1.501882e-05, 
    -1.501882e-05, -0.0001104672, -0.0002690957, -1.519242e-05, 4.069061e-06,
  -4.069061e-06, 1.519242e-05, 0.0002690957, 0.0001104672, 1.501882e-05, 
    1.501882e-05, 0.0001104672, 0.0002690957, 1.519242e-05, -4.069061e-06,
  -3.613859e-06, 1.373546e-05, 0.000883024, 0.0006720317, 0.0003086543, 
    0.0003086543, 0.0006720317, 0.000883024, 1.373546e-05, -3.613859e-06,
  0, -8.185861e-06, 0.001324375, 0.001488222, 0.001518787, 0.001518787, 
    0.001488222, 0.001324375, -8.185861e-06, 0,
  0, 0, 4.47583e-05, 0.0003188381, 0.0005194148, 0.0005194148, 0.0003188381, 
    4.47583e-05, 0, 0,
  0, 0, 0, -8.544845e-05, -0.0001391938, -0.0001391938, -8.544845e-05, 0, 0, 0,
  0, 0, 0, 5.822006e-09, 7.003699e-09, 7.003699e-09, 5.822006e-09, 0, 0, 0,
  0, 0, -1.331484e-08, -2.387134e-08, -2.873023e-08, -2.873023e-08, 
    -2.387134e-08, -1.331484e-08, 0, 0,
  0, -1.156787e-08, -2.344673e-08, -2.44924e-08, -2.523416e-08, 
    -2.523416e-08, -2.44924e-08, -2.344673e-08, -1.156787e-08, 0,
  5.861484e-10, -4.258139e-09, -1.553574e-08, -1.537197e-08, -1.533583e-08, 
    -1.533583e-08, -1.537197e-08, -1.553574e-08, -4.258139e-09, 5.861484e-10,
  3.122964e-10, -1.098778e-09, -4.864146e-09, -5.10307e-09, -5.883404e-09, 
    -5.883404e-09, -5.10307e-09, -4.864146e-09, -1.098778e-09, 3.122964e-10,
  -3.122964e-10, 1.098778e-09, 4.864146e-09, 5.10307e-09, 5.883404e-09, 
    5.883404e-09, 5.10307e-09, 4.864146e-09, 1.098778e-09, -3.122964e-10,
  -5.861484e-10, 4.258139e-09, 1.553574e-08, 1.537197e-08, 1.533583e-08, 
    1.533583e-08, 1.537197e-08, 1.553574e-08, 4.258139e-09, -5.861484e-10,
  0, 1.156787e-08, 2.344673e-08, 2.44924e-08, 2.523416e-08, 2.523416e-08, 
    2.44924e-08, 2.344673e-08, 1.156787e-08, 0,
  0, 0, 1.331484e-08, 2.387134e-08, 2.873023e-08, 2.873023e-08, 2.387134e-08, 
    1.331484e-08, 0, 0,
  0, 0, 0, -5.822006e-09, -7.003699e-09, -7.003699e-09, -5.822006e-09, 0, 0, 0,
  0, 0, 0, 0.0006145203, 0.0009423745, 0.0009423745, 0.0006145203, 0, 0, 0,
  0, 0, -0.000761056, -0.002291939, -0.003524209, -0.003524209, -0.002291939, 
    -0.000761056, 0, 0,
  0, -0.0002989912, -0.008313667, -0.009221511, -0.009451356, -0.009451356, 
    -0.009221511, -0.008313667, -0.0002989912, 0,
  3.446963e-05, -0.0001408909, -0.005538933, -0.004532514, -0.002400297, 
    -0.002400297, -0.004532514, -0.005538933, -0.0001408909, 3.446963e-05,
  2.833646e-05, -0.0001062195, -0.001694023, -0.0008527749, -0.0001504265, 
    -0.0001504265, -0.0008527749, -0.001694023, -0.0001062195, 2.833646e-05,
  -2.833646e-05, 0.0001062195, 0.001694023, 0.0008527749, 0.0001504265, 
    0.0001504265, 0.0008527749, 0.001694023, 0.0001062195, -2.833646e-05,
  -3.446963e-05, 0.0001408909, 0.005538933, 0.004532514, 0.002400297, 
    0.002400297, 0.004532514, 0.005538933, 0.0001408909, -3.446963e-05,
  0, 0.0002989912, 0.008313667, 0.009221511, 0.009451356, 0.009451356, 
    0.009221511, 0.008313667, 0.0002989912, 0,
  0, 0, 0.000761056, 0.002291939, 0.003524209, 0.003524209, 0.002291939, 
    0.000761056, 0, 0,
  0, 0, 0, -0.0006145203, -0.0009423745, -0.0009423745, -0.0006145203, 0, 0, 0,
  0, 0, 0, 0.0006018683, 0.0009309254, 0.0009309254, 0.0006018683, 0, 0, 0,
  0, 0, -0.0006946157, -0.002244339, -0.003476808, -0.003476808, 
    -0.002244339, -0.0006946157, 0, 0,
  0, -0.0002554863, -0.008243145, -0.009120974, -0.009326496, -0.009326496, 
    -0.009120974, -0.008243145, -0.0002554863, 0,
  3.265457e-05, -0.0001338267, -0.005477678, -0.004456076, -0.002324953, 
    -0.002324953, -0.004456076, -0.005477678, -0.0001338267, 3.265457e-05,
  2.809974e-05, -0.0001052244, -0.001671177, -0.0008233186, -0.0001416827, 
    -0.0001416827, -0.0008233186, -0.001671177, -0.0001052244, 2.809974e-05,
  -2.809974e-05, 0.0001052244, 0.001671177, 0.0008233186, 0.0001416827, 
    0.0001416827, 0.0008233186, 0.001671177, 0.0001052244, -2.809974e-05,
  -3.265457e-05, 0.0001338267, 0.005477678, 0.004456076, 0.002324953, 
    0.002324953, 0.004456076, 0.005477678, 0.0001338267, -3.265457e-05,
  0, 0.0002554863, 0.008243145, 0.009120974, 0.009326496, 0.009326496, 
    0.009120974, 0.008243145, 0.0002554863, 0,
  0, 0, 0.0006946157, 0.002244339, 0.003476808, 0.003476808, 0.002244339, 
    0.0006946157, 0, 0,
  0, 0, 0, -0.0006018683, -0.0009309254, -0.0009309254, -0.0006018683, 0, 0, 0,
  0, 0, 0, 0.000569397, 0.0008949178, 0.0008949178, 0.000569397, 0, 0, 0,
  0, 0, -0.0005744161, -0.002123483, -0.003339963, -0.003339963, 
    -0.002123483, -0.0005744161, 0, 0,
  0, -0.0001762706, -0.007975801, -0.008808539, -0.008962623, -0.008962623, 
    -0.008808539, -0.007975801, -0.0001762706, 0,
  2.965407e-05, -0.0001208219, -0.005282386, -0.004224174, -0.002135323, 
    -0.002135323, -0.004224174, -0.005282386, -0.0001208219, 2.965407e-05,
  2.726686e-05, -0.0001019677, -0.001603614, -0.0007551908, -0.0001242063, 
    -0.0001242063, -0.0007551908, -0.001603614, -0.0001019677, 2.726686e-05,
  -2.726686e-05, 0.0001019677, 0.001603614, 0.0007551908, 0.0001242063, 
    0.0001242063, 0.0007551908, 0.001603614, 0.0001019677, -2.726686e-05,
  -2.965407e-05, 0.0001208219, 0.005282386, 0.004224174, 0.002135323, 
    0.002135323, 0.004224174, 0.005282386, 0.0001208219, -2.965407e-05,
  0, 0.0001762706, 0.007975801, 0.008808539, 0.008962623, 0.008962623, 
    0.008808539, 0.007975801, 0.0001762706, 0,
  0, 0, 0.0005744161, 0.002123483, 0.003339963, 0.003339963, 0.002123483, 
    0.0005744161, 0, 0,
  0, 0, 0, -0.000569397, -0.0008949178, -0.0008949178, -0.000569397, 0, 0, 0,
  0, 0, 0, 0.0005155338, 0.0008197739, 0.0008197739, 0.0005155338, 0, 0, 0,
  0, 0, -0.0004545368, -0.001922653, -0.003058663, -0.003058663, 
    -0.001922653, -0.0004545368, 0, 0,
  0, -0.0001073958, -0.007372889, -0.008155355, -0.008276966, -0.008276966, 
    -0.008155355, -0.007372889, -0.0001073958, 0,
  2.58518e-05, -0.0001042298, -0.00488117, -0.003846478, -0.001887635, 
    -0.001887635, -0.003846478, -0.00488117, -0.0001042298, 2.58518e-05,
  2.493356e-05, -9.322522e-05, -0.001478728, -0.0006677705, -0.000103518, 
    -0.000103518, -0.0006677705, -0.001478728, -9.322522e-05, 2.493356e-05,
  -2.493356e-05, 9.322522e-05, 0.001478728, 0.0006677705, 0.000103518, 
    0.000103518, 0.0006677705, 0.001478728, 9.322522e-05, -2.493356e-05,
  -2.58518e-05, 0.0001042298, 0.00488117, 0.003846478, 0.001887635, 
    0.001887635, 0.003846478, 0.00488117, 0.0001042298, -2.58518e-05,
  0, 0.0001073958, 0.007372889, 0.008155355, 0.008276966, 0.008276966, 
    0.008155355, 0.007372889, 0.0001073958, 0,
  0, 0, 0.0004545368, 0.001922653, 0.003058663, 0.003058663, 0.001922653, 
    0.0004545368, 0, 0,
  0, 0, 0, -0.0005155338, -0.0008197739, -0.0008197739, -0.0005155338, 0, 0, 0,
  0, 0, 0, 0.0004427115, 0.0007094275, 0.0007094275, 0.0004427115, 0, 0, 0,
  0, 0, -0.0003462129, -0.001651167, -0.002646727, -0.002646727, 
    -0.001651167, -0.0003462129, 0, 0,
  0, -5.649689e-05, -0.006446572, -0.007149083, -0.007253477, -0.007253477, 
    -0.007149083, -0.006446572, -5.649689e-05, 0,
  2.146614e-05, -8.555062e-05, -0.004270537, -0.003329981, -0.001600625, 
    -0.001600625, -0.003329981, -0.004270537, -8.555062e-05, 2.146614e-05,
  2.142994e-05, -8.012012e-05, -0.00129395, -0.0005673318, -8.340323e-05, 
    -8.340323e-05, -0.0005673318, -0.00129395, -8.012012e-05, 2.142994e-05,
  -2.142994e-05, 8.012012e-05, 0.00129395, 0.0005673318, 8.340323e-05, 
    8.340323e-05, 0.0005673318, 0.00129395, 8.012012e-05, -2.142994e-05,
  -2.146614e-05, 8.555062e-05, 0.004270537, 0.003329981, 0.001600625, 
    0.001600625, 0.003329981, 0.004270537, 8.555062e-05, -2.146614e-05,
  0, 5.649689e-05, 0.006446572, 0.007149083, 0.007253477, 0.007253477, 
    0.007149083, 0.006446572, 5.649689e-05, 0,
  0, 0, 0.0003462129, 0.001651167, 0.002646727, 0.002646727, 0.001651167, 
    0.0003462129, 0, 0,
  0, 0, 0, -0.0004427115, -0.0007094275, -0.0007094275, -0.0004427115, 0, 0, 0,
  0, 0, 0, 0.0003578071, 0.0005763965, 0.0005763965, 0.0003578071, 0, 0, 0,
  0, 0, -0.0002518299, -0.001334621, -0.002150422, -0.002150422, 
    -0.001334621, -0.0002518299, 0, 0,
  0, -2.242266e-05, -0.005292843, -0.005883555, -0.005972451, -0.005972451, 
    -0.005883555, -0.005292843, -2.242266e-05, 0,
  1.685587e-05, -6.639662e-05, -0.003508329, -0.002713289, -0.001286073, 
    -0.001286073, -0.002713289, -0.003508329, -6.639662e-05, 1.685587e-05,
  1.727621e-05, -6.457946e-05, -0.001063868, -0.0004570856, -6.48932e-05, 
    -6.48932e-05, -0.0004570856, -0.001063868, -6.457946e-05, 1.727621e-05,
  -1.727621e-05, 6.457946e-05, 0.001063868, 0.0004570856, 6.48932e-05, 
    6.48932e-05, 0.0004570856, 0.001063868, 6.457946e-05, -1.727621e-05,
  -1.685587e-05, 6.639662e-05, 0.003508329, 0.002713289, 0.001286073, 
    0.001286073, 0.002713289, 0.003508329, 6.639662e-05, -1.685587e-05,
  0, 2.242266e-05, 0.005292843, 0.005883555, 0.005972451, 0.005972451, 
    0.005883555, 0.005292843, 2.242266e-05, 0,
  0, 0, 0.0002518299, 0.001334621, 0.002150422, 0.002150422, 0.001334621, 
    0.0002518299, 0, 0,
  0, 0, 0, -0.0003578071, -0.0005763965, -0.0005763965, -0.0003578071, 0, 0, 0,
  0, 0, 0, 0.0002673276, 0.0004321113, 0.0004321113, 0.0002673276, 0, 0, 0,
  0, 0, -0.0001719668, -0.0009972363, -0.001612196, -0.001612196, 
    -0.0009972363, -0.0001719668, 0, 0,
  0, -2.790395e-06, -0.004010062, -0.004465958, -0.004536331, -0.004536331, 
    -0.004465958, -0.004010062, -2.790395e-06, 0,
  1.229173e-05, -4.78558e-05, -0.002658849, -0.002041946, -0.0009582682, 
    -0.0009582682, -0.002041946, -0.002658849, -4.78558e-05, 1.229173e-05,
  1.285302e-05, -4.803204e-05, -0.0008069191, -0.0003415819, -4.758104e-05, 
    -4.758104e-05, -0.0003415819, -0.0008069191, -4.803204e-05, 1.285302e-05,
  -1.285302e-05, 4.803204e-05, 0.0008069191, 0.0003415819, 4.758104e-05, 
    4.758104e-05, 0.0003415819, 0.0008069191, 4.803204e-05, -1.285302e-05,
  -1.229173e-05, 4.78558e-05, 0.002658849, 0.002041946, 0.0009582682, 
    0.0009582682, 0.002041946, 0.002658849, 4.78558e-05, -1.229173e-05,
  0, 2.790395e-06, 0.004010062, 0.004465958, 0.004536331, 0.004536331, 
    0.004465958, 0.004010062, 2.790395e-06, 0,
  0, 0, 0.0001719668, 0.0009972363, 0.001612196, 0.001612196, 0.0009972363, 
    0.0001719668, 0, 0,
  0, 0, 0, -0.0002673276, -0.0004321113, -0.0004321113, -0.0002673276, 0, 0, 0,
  0, 0, 0, 0.0001758832, 0.0002848972, 0.0002848972, 0.0001758832, 0, 0, 0,
  0, 0, -0.0001047961, -0.0006561888, -0.001063018, -0.001063018, 
    -0.0006561888, -0.0001047961, 0, 0,
  0, 5.767954e-06, -0.002672944, -0.002982057, -0.003031253, -0.003031253, 
    -0.002982057, -0.002672944, 5.767954e-06, 0,
  7.908131e-06, -3.042558e-05, -0.001772953, -0.00135321, -0.0006300837, 
    -0.0006300837, -0.00135321, -0.001772953, -3.042558e-05, 7.908131e-06,
  8.413174e-06, -3.142826e-05, -0.000538476, -0.0002252401, -3.111303e-05, 
    -3.111303e-05, -0.0002252401, -0.000538476, -3.142826e-05, 8.413174e-06,
  -8.413174e-06, 3.142826e-05, 0.000538476, 0.0002252401, 3.111303e-05, 
    3.111303e-05, 0.0002252401, 0.000538476, 3.142826e-05, -8.413174e-06,
  -7.908131e-06, 3.042558e-05, 0.001772953, 0.00135321, 0.0006300837, 
    0.0006300837, 0.00135321, 0.001772953, 3.042558e-05, -7.908131e-06,
  0, -5.767954e-06, 0.002672944, 0.002982057, 0.003031253, 0.003031253, 
    0.002982057, 0.002672944, -5.767954e-06, 0,
  0, 0, 0.0001047961, 0.0006561888, 0.001063018, 0.001063018, 0.0006561888, 
    0.0001047961, 0, 0,
  0, 0, 0, -0.0001758832, -0.0002848972, -0.0002848972, -0.0001758832, 0, 0, 0,
  0, 0, 0, 8.623255e-05, 0.0001399608, 0.0001399608, 8.623255e-05, 0, 0, 0,
  0, 0, -4.760958e-05, -0.000321763, -0.0005222771, -0.0005222771, 
    -0.000321763, -4.760958e-05, 0, 0,
  0, 6.41051e-06, -0.001328308, -0.001486439, -0.001513435, -0.001513435, 
    -0.001486439, -0.001328308, 6.41051e-06, 0,
  3.767081e-06, -1.430753e-05, -0.0008826931, -0.0006711513, -0.0003103066, 
    -0.0003103066, -0.0006711513, -0.0008826931, -1.430753e-05, 3.767081e-06,
  4.104208e-06, -1.532345e-05, -0.000268516, -0.0001111782, -1.533146e-05, 
    -1.533146e-05, -0.0001111782, -0.000268516, -1.532345e-05, 4.104208e-06,
  -4.104208e-06, 1.532345e-05, 0.000268516, 0.0001111782, 1.533146e-05, 
    1.533146e-05, 0.0001111782, 0.000268516, 1.532345e-05, -4.104208e-06,
  -3.767081e-06, 1.430753e-05, 0.0008826931, 0.0006711513, 0.0003103066, 
    0.0003103066, 0.0006711513, 0.0008826931, 1.430753e-05, -3.767081e-06,
  0, -6.41051e-06, 0.001328308, 0.001486439, 0.001513435, 0.001513435, 
    0.001486439, 0.001328308, -6.41051e-06, 0,
  0, 0, 4.760958e-05, 0.000321763, 0.0005222771, 0.0005222771, 0.000321763, 
    4.760958e-05, 0, 0,
  0, 0, 0, -8.623255e-05, -0.0001399608, -0.0001399608, -8.623255e-05, 0, 0, 0,
  0, 0, 0, 5.82523e-09, 7.004086e-09, 7.004086e-09, 5.82523e-09, 0, 0, 0,
  0, 0, -1.334284e-08, -2.390036e-08, -2.875323e-08, -2.875323e-08, 
    -2.390036e-08, -1.334284e-08, 0, 0,
  0, -1.158092e-08, -2.343999e-08, -2.44425e-08, -2.516461e-08, 
    -2.516461e-08, -2.44425e-08, -2.343999e-08, -1.158092e-08, 0,
  5.863201e-10, -4.263859e-09, -1.552301e-08, -1.535468e-08, -1.534258e-08, 
    -1.534258e-08, -1.535468e-08, -1.552301e-08, -4.263859e-09, 5.863201e-10,
  3.123937e-10, -1.099315e-09, -4.861426e-09, -5.105515e-09, -5.903839e-09, 
    -5.903839e-09, -5.105515e-09, -4.861426e-09, -1.099315e-09, 3.123937e-10,
  -3.123937e-10, 1.099315e-09, 4.861426e-09, 5.105515e-09, 5.903839e-09, 
    5.903839e-09, 5.105515e-09, 4.861426e-09, 1.099315e-09, -3.123937e-10,
  -5.863201e-10, 4.263859e-09, 1.552301e-08, 1.535468e-08, 1.534258e-08, 
    1.534258e-08, 1.535468e-08, 1.552301e-08, 4.263859e-09, -5.863201e-10,
  0, 1.158092e-08, 2.343999e-08, 2.44425e-08, 2.516461e-08, 2.516461e-08, 
    2.44425e-08, 2.343999e-08, 1.158092e-08, 0,
  0, 0, 1.334284e-08, 2.390036e-08, 2.875323e-08, 2.875323e-08, 2.390036e-08, 
    1.334284e-08, 0, 0,
  0, 0, 0, -5.82523e-09, -7.004086e-09, -7.004086e-09, -5.82523e-09, 0, 0, 0,
  0, 0, 0, 0.0005071253, 0.0009713179, 0.0009713179, 0.0005071253, 0, 0, 0,
  0, -0.000122941, 0.0005770404, -0.001891851, -0.003632271, -0.003632271, 
    -0.001891851, 0.0005770404, -0.000122941, 0,
  0, 0.0005033952, -0.002340529, -0.008948468, -0.00943802, -0.00943802, 
    -0.008948468, -0.002340529, 0.0005033952, 0,
  4.86494e-05, -0.0001888947, -0.005456394, -0.004253624, -0.002438161, 
    -0.002438161, -0.004253624, -0.005456394, -0.0001888947, 4.86494e-05,
  2.325717e-05, -8.905558e-05, -0.001691033, -0.0008928971, -0.0001476524, 
    -0.0001476524, -0.0008928971, -0.001691033, -8.905558e-05, 2.325717e-05,
  -2.325717e-05, 8.905558e-05, 0.001691033, 0.0008928971, 0.0001476524, 
    0.0001476524, 0.0008928971, 0.001691033, 8.905558e-05, -2.325717e-05,
  -4.86494e-05, 0.0001888947, 0.005456394, 0.004253624, 0.002438161, 
    0.002438161, 0.004253624, 0.005456394, 0.0001888947, -4.86494e-05,
  0, -0.0005033952, 0.002340529, 0.008948468, 0.00943802, 0.00943802, 
    0.008948468, 0.002340529, -0.0005033952, 0,
  0, 0.000122941, -0.0005770404, 0.001891851, 0.003632271, 0.003632271, 
    0.001891851, -0.0005770404, 0.000122941, 0,
  0, 0, 0, -0.0005071253, -0.0009713179, -0.0009713179, -0.0005071253, 0, 0, 0,
  0, 0, 0, 0.000493344, 0.0009601261, 0.0009601261, 0.000493344, 0, 0, 0,
  0, -0.0001251832, 0.0005752536, -0.001841575, -0.003585364, -0.003585364, 
    -0.001841575, 0.0005752536, -0.0001251832, 0,
  0, 0.0005016397, -0.002295947, -0.008847, -0.00931478, -0.00931478, 
    -0.008847, -0.002295947, 0.0005016397, 0,
  4.504287e-05, -0.0001763244, -0.005395042, -0.004195032, -0.002360326, 
    -0.002360326, -0.004195032, -0.005395042, -0.0001763244, 4.504287e-05,
  2.358981e-05, -8.975093e-05, -0.001668034, -0.0008596442, -0.0001393442, 
    -0.0001393442, -0.0008596442, -0.001668034, -8.975093e-05, 2.358981e-05,
  -2.358981e-05, 8.975093e-05, 0.001668034, 0.0008596442, 0.0001393442, 
    0.0001393442, 0.0008596442, 0.001668034, 8.975093e-05, -2.358981e-05,
  -4.504287e-05, 0.0001763244, 0.005395042, 0.004195032, 0.002360326, 
    0.002360326, 0.004195032, 0.005395042, 0.0001763244, -4.504287e-05,
  0, -0.0005016397, 0.002295947, 0.008847, 0.00931478, 0.00931478, 0.008847, 
    0.002295947, -0.0005016397, 0,
  0, 0.0001251832, -0.0005752536, 0.001841575, 0.003585364, 0.003585364, 
    0.001841575, -0.0005752536, 0.0001251832, 0,
  0, 0, 0, -0.000493344, -0.0009601261, -0.0009601261, -0.000493344, 0, 0, 0,
  0, 0, 0, 0.0004607817, 0.000924008, 0.000924008, 0.0004607817, 0, 0, 0,
  0, -0.0001248465, 0.0005574753, -0.001720755, -0.003447955, -0.003447955, 
    -0.001720755, 0.0005574753, -0.0001248465, 0,
  0, 0.0004885047, -0.002183635, -0.00853559, -0.008954303, -0.008954303, 
    -0.00853559, -0.002183635, 0.0004885047, 0,
  3.923894e-05, -0.0001540941, -0.005204882, -0.003996574, -0.00216685, 
    -0.00216685, -0.003996574, -0.005204882, -0.0001540941, 3.923894e-05,
  2.362618e-05, -8.927784e-05, -0.001599355, -0.0007861073, -0.0001223268, 
    -0.0001223268, -0.0007861073, -0.001599355, -8.927784e-05, 2.362618e-05,
  -2.362618e-05, 8.927784e-05, 0.001599355, 0.0007861073, 0.0001223268, 
    0.0001223268, 0.0007861073, 0.001599355, 8.927784e-05, -2.362618e-05,
  -3.923894e-05, 0.0001540941, 0.005204882, 0.003996574, 0.00216685, 
    0.00216685, 0.003996574, 0.005204882, 0.0001540941, -3.923894e-05,
  0, -0.0004885047, 0.002183635, 0.00853559, 0.008954303, 0.008954303, 
    0.00853559, 0.002183635, -0.0004885047, 0,
  0, 0.0001248465, -0.0005574753, 0.001720755, 0.003447955, 0.003447955, 
    0.001720755, -0.0005574753, 0.0001248465, 0,
  0, 0, 0, -0.0004607817, -0.000924008, -0.000924008, -0.0004607817, 0, 0, 0,
  0, 0, 0, 0.0004127499, 0.0008472838, 0.0008472838, 0.0004127499, 0, 0, 0,
  0, -0.0001174738, 0.000513422, -0.001541335, -0.003160817, -0.003160817, 
    -0.001541335, 0.000513422, -0.0001174738, 0,
  0, 0.0004535116, -0.001988313, -0.007900783, -0.00827109, -0.00827109, 
    -0.007900783, -0.001988313, 0.0004535116, 0,
  3.298846e-05, -0.0001292149, -0.004817074, -0.003653675, -0.001915359, 
    -0.001915359, -0.003653675, -0.004817074, -0.0001292149, 3.298846e-05,
  2.209667e-05, -8.322528e-05, -0.001472444, -0.0006939937, -0.0001019367, 
    -0.0001019367, -0.0006939937, -0.001472444, -8.322528e-05, 2.209667e-05,
  -2.209667e-05, 8.322528e-05, 0.001472444, 0.0006939937, 0.0001019367, 
    0.0001019367, 0.0006939937, 0.001472444, 8.322528e-05, -2.209667e-05,
  -3.298846e-05, 0.0001292149, 0.004817074, 0.003653675, 0.001915359, 
    0.001915359, 0.003653675, 0.004817074, 0.0001292149, -3.298846e-05,
  0, -0.0004535116, 0.001988313, 0.007900783, 0.00827109, 0.00827109, 
    0.007900783, 0.001988313, -0.0004535116, 0,
  0, 0.0001174738, -0.000513422, 0.001541335, 0.003160817, 0.003160817, 
    0.001541335, -0.000513422, 0.0001174738, 0,
  0, 0, 0, -0.0004127499, -0.0008472838, -0.0008472838, -0.0004127499, 0, 0, 0,
  0, 0, 0, 0.000351859, 0.0007338061, 0.0007338061, 0.000351859, 0, 0, 0,
  0, -0.0001035608, 0.0004460113, -0.001313798, -0.002737319, -0.002737319, 
    -0.001313798, 0.0004460113, -0.0001035608, 0,
  0, 0.0003970476, -0.001716495, -0.006928134, -0.007249506, -0.007249506, 
    -0.006928134, -0.001716495, 0.0003970476, 0,
  2.664342e-05, -0.0001038137, -0.004223715, -0.003172668, -0.00162399, 
    -0.00162399, -0.003172668, -0.004223715, -0.0001038137, 2.664342e-05,
  1.928389e-05, -7.248516e-05, -0.001285968, -0.0005888975, -8.213058e-05, 
    -8.213058e-05, -0.0005888975, -0.001285968, -7.248516e-05, 1.928389e-05,
  -1.928389e-05, 7.248516e-05, 0.001285968, 0.0005888975, 8.213058e-05, 
    8.213058e-05, 0.0005888975, 0.001285968, 7.248516e-05, -1.928389e-05,
  -2.664342e-05, 0.0001038137, 0.004223715, 0.003172668, 0.00162399, 
    0.00162399, 0.003172668, 0.004223715, 0.0001038137, -2.664342e-05,
  0, -0.0003970476, 0.001716495, 0.006928134, 0.007249506, 0.007249506, 
    0.006928134, 0.001716495, -0.0003970476, 0,
  0, 0.0001035608, -0.0004460113, 0.001313798, 0.002737319, 0.002737319, 
    0.001313798, -0.0004460113, 0.0001035608, 0,
  0, 0, 0, -0.000351859, -0.0007338061, -0.0007338061, -0.000351859, 0, 0, 0,
  0, 0, 0, 0.0002829162, 0.0005965838, 0.0005965838, 0.0002829162, 0, 0, 0,
  0, -8.528172e-05, 0.0003635667, -0.001056253, -0.0022255, -0.0022255, 
    -0.001056253, 0.0003635667, -8.528172e-05, 0,
  0, 0.0003256902, -0.001394031, -0.005705225, -0.005970362, -0.005970362, 
    -0.005705225, -0.001394031, 0.0003256902, 0,
  2.044338e-05, -7.914679e-05, -0.00347805, -0.002591366, -0.001304716, 
    -0.001304716, -0.002591366, -0.00347805, -7.914679e-05, 2.044338e-05,
  1.572823e-05, -5.902622e-05, -0.001055357, -0.000473982, -6.393938e-05, 
    -6.393938e-05, -0.000473982, -0.001055357, -5.902622e-05, 1.572823e-05,
  -1.572823e-05, 5.902622e-05, 0.001055357, 0.000473982, 6.393938e-05, 
    6.393938e-05, 0.000473982, 0.001055357, 5.902622e-05, -1.572823e-05,
  -2.044338e-05, 7.914679e-05, 0.00347805, 0.002591366, 0.001304716, 
    0.001304716, 0.002591366, 0.00347805, 7.914679e-05, -2.044338e-05,
  0, -0.0003256902, 0.001394031, 0.005705225, 0.005970362, 0.005970362, 
    0.005705225, 0.001394031, -0.0003256902, 0,
  0, 8.528172e-05, -0.0003635667, 0.001056253, 0.0022255, 0.0022255, 
    0.001056253, -0.0003635667, 8.528172e-05, 0,
  0, 0, 0, -0.0002829162, -0.0005965838, -0.0005965838, -0.0002829162, 0, 0, 0,
  0, 0, 0, 0.0002105939, 0.000447504, 0.000447504, 0.0002105939, 0, 0, 0,
  0, -6.459056e-05, 0.0002734499, -0.0007861596, -0.001669488, -0.001669488, 
    -0.0007861596, 0.0002734499, -6.459056e-05, 0,
  0, 0.0002460892, -0.001046096, -0.004334302, -0.004536202, -0.004536202, 
    -0.004334302, -0.001046096, 0.0002460892, 0,
  1.460284e-05, -5.613481e-05, -0.002642252, -0.001954187, -0.0009721543, 
    -0.0009721543, -0.001954187, -0.002642252, -5.613481e-05, 1.460284e-05,
  1.181465e-05, -4.427704e-05, -0.0007992044, -0.0003539496, -4.692788e-05, 
    -4.692788e-05, -0.0003539496, -0.0007992044, -4.427704e-05, 1.181465e-05,
  -1.181465e-05, 4.427704e-05, 0.0007992044, 0.0003539496, 4.692788e-05, 
    4.692788e-05, 0.0003539496, 0.0007992044, 4.427704e-05, -1.181465e-05,
  -1.460284e-05, 5.613481e-05, 0.002642252, 0.001954187, 0.0009721543, 
    0.0009721543, 0.001954187, 0.002642252, 5.613481e-05, -1.460284e-05,
  0, -0.0002460892, 0.001046096, 0.004334302, 0.004536202, 0.004536202, 
    0.004334302, 0.001046096, -0.0002460892, 0,
  0, 6.459056e-05, -0.0002734499, 0.0007861596, 0.001669488, 0.001669488, 
    0.0007861596, -0.0002734499, 6.459056e-05, 0,
  0, 0, 0, -0.0002105939, -0.000447504, -0.000447504, -0.0002105939, 0, 0, 0,
  0, 0, 0, 0.0001381627, 0.0002952171, 0.0002952171, 0.0001381627, 0, 0, 0,
  0, -4.292298e-05, 0.0001808726, -0.0005157209, -0.00110146, -0.00110146, 
    -0.0005157209, 0.0001808726, -4.292298e-05, 0,
  0, 0.0001632886, -0.0006909294, -0.00289724, -0.003032865, -0.003032865, 
    -0.00289724, -0.0006909294, 0.0001632886, 0,
  9.211845e-06, -3.513769e-05, -0.00176618, -0.001297592, -0.0006393747, 
    -0.0006393747, -0.001297592, -0.00176618, -3.513769e-05, 9.211845e-06,
  7.80042e-06, -2.919402e-05, -0.0005327126, -0.0002333162, -3.072609e-05, 
    -3.072609e-05, -0.0002333162, -0.0005327126, -2.919402e-05, 7.80042e-06,
  -7.80042e-06, 2.919402e-05, 0.0005327126, 0.0002333162, 3.072609e-05, 
    3.072609e-05, 0.0002333162, 0.0005327126, 2.919402e-05, -7.80042e-06,
  -9.211845e-06, 3.513769e-05, 0.00176618, 0.001297592, 0.0006393747, 
    0.0006393747, 0.001297592, 0.00176618, 3.513769e-05, -9.211845e-06,
  0, -0.0001632886, 0.0006909294, 0.00289724, 0.003032865, 0.003032865, 
    0.00289724, 0.0006909294, -0.0001632886, 0,
  0, 4.292298e-05, -0.0001808726, 0.0005157209, 0.00110146, 0.00110146, 
    0.0005157209, -0.0001808726, 4.292298e-05, 0,
  0, 0, 0, -0.0001381627, -0.0002952171, -0.0002952171, -0.0001381627, 0, 0, 0,
  0, 0, 0, 6.754683e-05, 0.0001451101, 0.0001451101, 6.754683e-05, 0, 0, 0,
  0, -2.121002e-05, 8.90798e-05, -0.0002521111, -0.0005414747, -0.0005414747, 
    -0.0002521111, 8.90798e-05, -2.121002e-05, 0,
  0, 8.059232e-05, -0.0003399263, -0.00144566, -0.001515442, -0.001515442, 
    -0.00144566, -0.0003399263, 8.059232e-05, 0,
  4.301308e-06, -1.626051e-05, -0.0008812804, -0.0006449149, -0.0003151101, 
    -0.0003151101, -0.0006449149, -0.0008812804, -1.626051e-05, 4.301308e-06,
  3.837732e-06, -1.434243e-05, -0.0002654715, -0.0001151896, -1.516404e-05, 
    -1.516404e-05, -0.0001151896, -0.0002654715, -1.434243e-05, 3.837732e-06,
  -3.837732e-06, 1.434243e-05, 0.0002654715, 0.0001151896, 1.516404e-05, 
    1.516404e-05, 0.0001151896, 0.0002654715, 1.434243e-05, -3.837732e-06,
  -4.301308e-06, 1.626051e-05, 0.0008812804, 0.0006449149, 0.0003151101, 
    0.0003151101, 0.0006449149, 0.0008812804, 1.626051e-05, -4.301308e-06,
  0, -8.059232e-05, 0.0003399263, 0.00144566, 0.001515442, 0.001515442, 
    0.00144566, 0.0003399263, -8.059232e-05, 0,
  0, 2.121002e-05, -8.90798e-05, 0.0002521111, 0.0005414747, 0.0005414747, 
    0.0002521111, -8.90798e-05, 2.121002e-05, 0,
  0, 0, 0, -6.754683e-05, -0.0001451101, -0.0001451101, -6.754683e-05, 0, 0, 0,
  0, 0, 0, 5.804671e-09, 7.008032e-09, 7.008032e-09, 5.804671e-09, 0, 0, 0,
  0, 2.319781e-09, -4.230289e-09, -2.381888e-08, -2.878978e-08, 
    -2.878978e-08, -2.381888e-08, -4.230289e-09, 2.319781e-09, 0,
  0, -4.599584e-09, -1.879162e-08, -2.450905e-08, -2.506749e-08, 
    -2.506749e-08, -2.450905e-08, -1.879162e-08, -4.599584e-09, 0,
  8.882792e-10, -4.862396e-09, -1.511646e-08, -1.50993e-08, -1.539255e-08, 
    -1.539255e-08, -1.50993e-08, -1.511646e-08, -4.862396e-09, 8.882792e-10,
  2.049165e-10, -9.173195e-10, -4.975775e-09, -5.1423e-09, -5.910174e-09, 
    -5.910174e-09, -5.1423e-09, -4.975775e-09, -9.173195e-10, 2.049165e-10,
  -2.049165e-10, 9.173195e-10, 4.975775e-09, 5.1423e-09, 5.910174e-09, 
    5.910174e-09, 5.1423e-09, 4.975775e-09, 9.173195e-10, -2.049165e-10,
  -8.882792e-10, 4.862396e-09, 1.511646e-08, 1.50993e-08, 1.539255e-08, 
    1.539255e-08, 1.50993e-08, 1.511646e-08, 4.862396e-09, -8.882792e-10,
  0, 4.599584e-09, 1.879162e-08, 2.450905e-08, 2.506749e-08, 2.506749e-08, 
    2.450905e-08, 1.879162e-08, 4.599584e-09, 0,
  0, -2.319781e-09, 4.230289e-09, 2.381888e-08, 2.878978e-08, 2.878978e-08, 
    2.381888e-08, 4.230289e-09, -2.319781e-09, 0,
  0, 0, 0, -5.804671e-09, -7.008032e-09, -7.008032e-09, -5.804671e-09, 0, 0, 0,
  0, 0, 0, 0.0005110904, 0.0009751136, 0.0009751136, 0.0005110904, 0, 0, 0,
  0, -0.0001232052, 0.0005791325, -0.0019067, -0.003646616, -0.003646616, 
    -0.0019067, 0.0005791325, -0.0001232052, 0,
  0, 0.0005050731, -0.002350952, -0.008924956, -0.009382538, -0.009382538, 
    -0.008924956, -0.002350952, 0.0005050731, 0,
  4.980121e-05, -0.0001931989, -0.005442988, -0.004234629, -0.002442166, 
    -0.002442166, -0.004234629, -0.005442988, -0.0001931989, 4.980121e-05,
  2.342554e-05, -8.968446e-05, -0.001682935, -0.0008943132, -0.0001501193, 
    -0.0001501193, -0.0008943132, -0.001682935, -8.968446e-05, 2.342554e-05,
  -2.342554e-05, 8.968446e-05, 0.001682935, 0.0008943132, 0.0001501193, 
    0.0001501193, 0.0008943132, 0.001682935, 8.968446e-05, -2.342554e-05,
  -4.980121e-05, 0.0001931989, 0.005442988, 0.004234629, 0.002442166, 
    0.002442166, 0.004234629, 0.005442988, 0.0001931989, -4.980121e-05,
  0, -0.0005050731, 0.002350952, 0.008924956, 0.009382538, 0.009382538, 
    0.008924956, 0.002350952, -0.0005050731, 0,
  0, 0.0001232052, -0.0005791325, 0.0019067, 0.003646616, 0.003646616, 
    0.0019067, -0.0005791325, 0.0001232052, 0,
  0, 0, 0, -0.0005110904, -0.0009751136, -0.0009751136, -0.0005110904, 0, 0, 0,
  0, 0, 0, 0.0004972908, 0.0009639504, 0.0009639504, 0.0004972908, 0, 0, 0,
  0, -0.0001254825, 0.0005774138, -0.001856323, -0.003599732, -0.003599732, 
    -0.001856323, 0.0005774138, -0.0001254825, 0,
  0, 0.0005033801, -0.002306366, -0.008823977, -0.009260577, -0.009260577, 
    -0.008823977, -0.002306366, 0.0005033801, 0,
  4.618923e-05, -0.0001806051, -0.005381955, -0.004176188, -0.002364439, 
    -0.002364439, -0.004176188, -0.005381955, -0.0001806051, 4.618923e-05,
  2.375904e-05, -9.038047e-05, -0.001660131, -0.0008612028, -0.0001416985, 
    -0.0001416985, -0.0008612028, -0.001660131, -9.038047e-05, 2.375904e-05,
  -2.375904e-05, 9.038047e-05, 0.001660131, 0.0008612028, 0.0001416985, 
    0.0001416985, 0.0008612028, 0.001660131, 9.038047e-05, -2.375904e-05,
  -4.618923e-05, 0.0001806051, 0.005381955, 0.004176188, 0.002364439, 
    0.002364439, 0.004176188, 0.005381955, 0.0001806051, -4.618923e-05,
  0, -0.0005033801, 0.002306366, 0.008823977, 0.009260577, 0.009260577, 
    0.008823977, 0.002306366, -0.0005033801, 0,
  0, 0.0001254825, -0.0005774138, 0.001856323, 0.003599732, 0.003599732, 
    0.001856323, -0.0005774138, 0.0001254825, 0,
  0, 0, 0, -0.0004972908, -0.0009639504, -0.0009639504, -0.0004972908, 0, 0, 0,
  0, 0, 0, 0.0004646453, 0.0009277874, 0.0009277874, 0.0004646453, 0, 0, 0,
  0, -0.0001251925, 0.0005597036, -0.001735174, -0.003462107, -0.003462107, 
    -0.001735174, 0.0005597036, -0.0001251925, 0,
  0, 0.0004903096, -0.002193888, -0.008513852, -0.008902945, -0.008902945, 
    -0.008513852, -0.002193888, 0.0004903096, 0,
  4.035887e-05, -0.0001582718, -0.005192575, -0.0039785, -0.002171342, 
    -0.002171342, -0.0039785, -0.005192575, -0.0001582718, 4.035887e-05,
  2.379059e-05, -8.98889e-05, -0.001591897, -0.0007879224, -0.0001243996, 
    -0.0001243996, -0.0007879224, -0.001591897, -8.98889e-05, 2.379059e-05,
  -2.379059e-05, 8.98889e-05, 0.001591897, 0.0007879224, 0.0001243996, 
    0.0001243996, 0.0007879224, 0.001591897, 8.98889e-05, -2.379059e-05,
  -4.035887e-05, 0.0001582718, 0.005192575, 0.0039785, 0.002171342, 
    0.002171342, 0.0039785, 0.005192575, 0.0001582718, -4.035887e-05,
  0, -0.0004903096, 0.002193888, 0.008513852, 0.008902945, 0.008902945, 
    0.008513852, 0.002193888, -0.0004903096, 0,
  0, 0.0001251925, -0.0005597036, 0.001735174, 0.003462107, 0.003462107, 
    0.001735174, -0.0005597036, 0.0001251925, 0,
  0, 0, 0, -0.0004646453, -0.0009277874, -0.0009277874, -0.0004646453, 0, 0, 0,
  0, 0, 0, 0.0004163565, 0.0008508377, 0.0008508377, 0.0004163565, 0, 0, 0,
  0, -0.0001178382, 0.0005156007, -0.001554788, -0.003174104, -0.003174104, 
    -0.001554788, 0.0005156007, -0.0001178382, 0,
  0, 0.0004552921, -0.001998015, -0.007881463, -0.008224366, -0.008224366, 
    -0.007881463, -0.001998015, 0.0004552921, 0,
  3.402655e-05, -0.0001330857, -0.004806186, -0.003637122, -0.001920068, 
    -0.001920068, -0.003637122, -0.004806186, -0.0001330857, 3.402655e-05,
  2.22479e-05, -8.378804e-05, -0.001465671, -0.0006959632, -0.0001036839, 
    -0.0001036839, -0.0006959632, -0.001465671, -8.378804e-05, 2.22479e-05,
  -2.22479e-05, 8.378804e-05, 0.001465671, 0.0006959632, 0.0001036839, 
    0.0001036839, 0.0006959632, 0.001465671, 8.378804e-05, -2.22479e-05,
  -3.402655e-05, 0.0001330857, 0.004806186, 0.003637122, 0.001920068, 
    0.001920068, 0.003637122, 0.004806186, 0.0001330857, -3.402655e-05,
  0, -0.0004552921, 0.001998015, 0.007881463, 0.008224366, 0.008224366, 
    0.007881463, 0.001998015, -0.0004552921, 0,
  0, 0.0001178382, -0.0005156007, 0.001554788, 0.003174104, 0.003174104, 
    0.001554788, -0.0005156007, 0.0001178382, 0,
  0, 0, 0, -0.0004163565, -0.0008508377, -0.0008508377, -0.0004163565, 0, 0, 0,
  0, 0, 0, 0.000355047, 0.0007369739, 0.0007369739, 0.000355047, 0, 0, 0,
  0, -0.0001039136, 0.000448019, -0.001325687, -0.002749153, -0.002749153, 
    -0.001325687, 0.000448019, -0.0001039136, 0,
  0, 0.0003987052, -0.001725244, -0.006912369, -0.007209442, -0.007209442, 
    -0.006912369, -0.001725244, 0.0003987052, 0,
  2.754993e-05, -0.0001071937, -0.004214888, -0.003158372, -0.001628536, 
    -0.001628536, -0.003158372, -0.004214888, -0.0001071937, 2.754993e-05,
  1.941581e-05, -7.297657e-05, -0.001280167, -0.000590838, -8.356683e-05, 
    -8.356683e-05, -0.000590838, -0.001280167, -7.297657e-05, 1.941581e-05,
  -1.941581e-05, 7.297657e-05, 0.001280167, 0.000590838, 8.356683e-05, 
    8.356683e-05, 0.000590838, 0.001280167, 7.297657e-05, -1.941581e-05,
  -2.754993e-05, 0.0001071937, 0.004214888, 0.003158372, 0.001628536, 
    0.001628536, 0.003158372, 0.004214888, 0.0001071937, -2.754993e-05,
  0, -0.0003987052, 0.001725244, 0.006912369, 0.007209442, 0.007209442, 
    0.006912369, 0.001725244, -0.0003987052, 0,
  0, 0.0001039136, -0.000448019, 0.001325687, 0.002749153, 0.002749153, 
    0.001325687, -0.000448019, 0.0001039136, 0,
  0, 0, 0, -0.000355047, -0.0007369739, -0.0007369739, -0.000355047, 0, 0, 0,
  0, 0, 0, 0.0002855763, 0.0005992496, 0.0005992496, 0.0002855763, 0, 0, 0,
  0, -8.559917e-05, 0.0003653085, -0.001066172, -0.002235452, -0.002235452, 
    -0.001066172, 0.0003653085, -8.559917e-05, 0,
  0, 0.000327143, -0.001401504, -0.005693769, -0.005938564, -0.005938564, 
    -0.005693769, -0.001401504, 0.000327143, 0,
  2.118585e-05, -8.191521e-05, -0.00347171, -0.002579907, -0.001308785, 
    -0.001308785, -0.002579907, -0.00347171, -8.191521e-05, 2.118585e-05,
  1.583643e-05, -5.942961e-05, -0.001050762, -0.0004757417, -6.508073e-05, 
    -6.508073e-05, -0.0004757417, -0.001050762, -5.942961e-05, 1.583643e-05,
  -1.583643e-05, 5.942961e-05, 0.001050762, 0.0004757417, 6.508073e-05, 
    6.508073e-05, 0.0004757417, 0.001050762, 5.942961e-05, -1.583643e-05,
  -2.118585e-05, 8.191521e-05, 0.00347171, 0.002579907, 0.001308785, 
    0.001308785, 0.002579907, 0.00347171, 8.191521e-05, -2.118585e-05,
  0, -0.000327143, 0.001401504, 0.005693769, 0.005938564, 0.005938564, 
    0.005693769, 0.001401504, -0.000327143, 0,
  0, 8.559917e-05, -0.0003653085, 0.001066172, 0.002235452, 0.002235452, 
    0.001066172, -0.0003653085, 8.559917e-05, 0,
  0, 0, 0, -0.0002855763, -0.0005992496, -0.0005992496, -0.0002855763, 0, 0, 0,
  0, 0, 0, 0.00021265, 0.000449594, 0.000449594, 0.00021265, 0, 0, 0,
  0, -6.485327e-05, 0.0002748477, -0.0007938269, -0.001677288, -0.001677288, 
    -0.0007938269, 0.0002748477, -6.485327e-05, 0,
  0, 0.0002472673, -0.00105202, -0.004327347, -0.004513612, -0.004513612, 
    -0.004327347, -0.00105202, 0.0002472673, 0,
  1.51612e-05, -5.821702e-05, -0.0026385, -0.001945966, -0.0009755426, 
    -0.0009755426, -0.001945966, -0.0026385, -5.821702e-05, 1.51612e-05,
  1.189718e-05, -4.458491e-05, -0.000795964, -0.0003554224, -4.778522e-05, 
    -4.778522e-05, -0.0003554224, -0.000795964, -4.458491e-05, 1.189718e-05,
  -1.189718e-05, 4.458491e-05, 0.000795964, 0.0003554224, 4.778522e-05, 
    4.778522e-05, 0.0003554224, 0.000795964, 4.458491e-05, -1.189718e-05,
  -1.51612e-05, 5.821702e-05, 0.0026385, 0.001945966, 0.0009755426, 
    0.0009755426, 0.001945966, 0.0026385, 5.821702e-05, -1.51612e-05,
  0, -0.0002472673, 0.00105202, 0.004327347, 0.004513612, 0.004513612, 
    0.004327347, 0.00105202, -0.0002472673, 0,
  0, 6.485327e-05, -0.0002748477, 0.0007938269, 0.001677288, 0.001677288, 
    0.0007938269, -0.0002748477, 6.485327e-05, 0,
  0, 0, 0, -0.00021265, -0.000449594, -0.000449594, -0.00021265, 0, 0, 0,
  0, 0, 0, 0.0001395506, 0.0002966736, 0.0002966736, 0.0001395506, 0, 0, 0,
  0, -4.311253e-05, 0.0001818528, -0.000520897, -0.001106895, -0.001106895, 
    -0.000520897, 0.0001818528, -4.311253e-05, 0,
  0, 0.0001641228, -0.0006950366, -0.002894199, -0.003019516, -0.003019516, 
    -0.002894199, -0.0006950366, 0.0001641228, 0,
  9.574579e-06, -3.649069e-05, -0.001764653, -0.001292788, -0.0006419583, 
    -0.0006419583, -0.001292788, -0.001764653, -3.649069e-05, 9.574579e-06,
  7.856769e-06, -2.940429e-05, -0.0005308443, -0.0002344245, -3.13057e-05, 
    -3.13057e-05, -0.0002344245, -0.0005308443, -2.940429e-05, 7.856769e-06,
  -7.856769e-06, 2.940429e-05, 0.0005308443, 0.0002344245, 3.13057e-05, 
    3.13057e-05, 0.0002344245, 0.0005308443, 2.940429e-05, -7.856769e-06,
  -9.574579e-06, 3.649069e-05, 0.001764653, 0.001292788, 0.0006419583, 
    0.0006419583, 0.001292788, 0.001764653, 3.649069e-05, -9.574579e-06,
  0, -0.0001641228, 0.0006950366, 0.002894199, 0.003019516, 0.003019516, 
    0.002894199, 0.0006950366, -0.0001641228, 0,
  0, 4.311253e-05, -0.0001818528, 0.000520897, 0.001106895, 0.001106895, 
    0.000520897, -0.0001818528, 4.311253e-05, 0,
  0, 0, 0, -0.0001395506, -0.0002966736, -0.0002966736, -0.0001395506, 0, 0, 0,
  0, 0, 0, 6.823079e-05, 0.0001458607, 0.0001458607, 6.823079e-05, 0, 0, 0,
  0, -2.130998e-05, 8.958419e-05, -0.0002546627, -0.0005442753, 
    -0.0005442753, -0.0002546627, 8.958419e-05, -2.130998e-05, 0,
  0, 8.10249e-05, -0.0003420194, -0.001444988, -0.001509905, -0.001509905, 
    -0.001444988, -0.0003420194, 8.10249e-05, 0,
  4.472497e-06, -1.689914e-05, -0.0008810312, -0.0006430848, -0.000316673, 
    -0.000316673, -0.0006430848, -0.0008810312, -1.689914e-05, 4.472497e-06,
  3.866233e-06, -1.444882e-05, -0.0002647389, -0.0001158388, -1.546205e-05, 
    -1.546205e-05, -0.0001158388, -0.0002647389, -1.444882e-05, 3.866233e-06,
  -3.866233e-06, 1.444882e-05, 0.0002647389, 0.0001158388, 1.546205e-05, 
    1.546205e-05, 0.0001158388, 0.0002647389, 1.444882e-05, -3.866233e-06,
  -4.472497e-06, 1.689914e-05, 0.0008810312, 0.0006430848, 0.000316673, 
    0.000316673, 0.0006430848, 0.0008810312, 1.689914e-05, -4.472497e-06,
  0, -8.10249e-05, 0.0003420194, 0.001444988, 0.001509905, 0.001509905, 
    0.001444988, 0.0003420194, -8.10249e-05, 0,
  0, 2.130998e-05, -8.958419e-05, 0.0002546627, 0.0005442753, 0.0005442753, 
    0.0002546627, -8.958419e-05, 2.130998e-05, 0,
  0, 0, 0, -6.823079e-05, -0.0001458607, -0.0001458607, -6.823079e-05, 0, 0, 0,
  0, 0, 0, 5.808406e-09, 7.008185e-09, 7.008185e-09, 5.808406e-09, 0, 0, 0,
  0, 2.323635e-09, -4.243433e-09, -2.384734e-08, -2.881204e-08, 
    -2.881204e-08, -2.384734e-08, -4.243433e-09, 2.323635e-09, 0,
  0, -4.609836e-09, -1.879897e-08, -2.446902e-08, -2.500002e-08, 
    -2.500002e-08, -2.446902e-08, -1.879897e-08, -4.609836e-09, 0,
  8.882624e-10, -4.868089e-09, -1.509725e-08, -1.507616e-08, -1.539884e-08, 
    -1.539884e-08, -1.507616e-08, -1.509725e-08, -4.868089e-09, 8.882624e-10,
  2.051505e-10, -9.183869e-10, -4.972821e-09, -5.141223e-09, -5.929314e-09, 
    -5.929314e-09, -5.141223e-09, -4.972821e-09, -9.183869e-10, 2.051505e-10,
  -2.051505e-10, 9.183869e-10, 4.972821e-09, 5.141223e-09, 5.929314e-09, 
    5.929314e-09, 5.141223e-09, 4.972821e-09, 9.183869e-10, -2.051505e-10,
  -8.882624e-10, 4.868089e-09, 1.509725e-08, 1.507616e-08, 1.539884e-08, 
    1.539884e-08, 1.507616e-08, 1.509725e-08, 4.868089e-09, -8.882624e-10,
  0, 4.609836e-09, 1.879897e-08, 2.446902e-08, 2.500002e-08, 2.500002e-08, 
    2.446902e-08, 1.879897e-08, 4.609836e-09, 0,
  0, -2.323635e-09, 4.243433e-09, 2.384734e-08, 2.881204e-08, 2.881204e-08, 
    2.384734e-08, 4.243433e-09, -2.323635e-09, 0,
  0, 0, 0, -5.808406e-09, -7.008185e-09, -7.008185e-09, -5.808406e-09, 0, 0, 0 ;
}
